-- p2_grms_qsys.vhd

-- Generated using ACDS version 13.0sp1 232 at 2023.01.05.16:32:28

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity p2_grms_qsys is
	port (
		clk_clk                              : in    std_logic                     := '0';             --                            clk.clk
		reset_reset_n                        : in    std_logic                     := '0';             --                          reset.reset_n
		pi_grms_external_connection_export   : out   std_logic_vector(3 downto 0);                     --    pi_grms_external_connection.export
		ph_grms_external_connection_export   : out   std_logic_vector(3 downto 0);                     --    ph_grms_external_connection.export
		pg_grms_external_connection_export   : out   std_logic_vector(6 downto 0);                     --    pg_grms_external_connection.export
		pf_grms_external_connection_export   : out   std_logic_vector(6 downto 0);                     --    pf_grms_external_connection.export
		pe_grms_external_connection_export   : out   std_logic_vector(7 downto 0);                     --    pe_grms_external_connection.export
		pd_grms_external_connection_export   : out   std_logic_vector(7 downto 0);                     --    pd_grms_external_connection.export
		pc_grms_external_connection_export   : out   std_logic;                                        --    pc_grms_external_connection.export
		pb_grms_external_connection_export   : in    std_logic_vector(3 downto 0)  := (others => '0'); --    pb_grms_external_connection.export
		pa_grms_external_connection_export   : in    std_logic_vector(7 downto 0)  := (others => '0'); --    pa_grms_external_connection.export
		lcd_16207_grms_external_RS           : out   std_logic;                                        --        lcd_16207_grms_external.RS
		lcd_16207_grms_external_RW           : out   std_logic;                                        --                               .RW
		lcd_16207_grms_external_data         : inout std_logic_vector(7 downto 0)  := (others => '0'); --                               .data
		lcd_16207_grms_external_E            : out   std_logic;                                        --                               .E
		new_sdram_controller_grms_wire_addr  : out   std_logic_vector(11 downto 0);                    -- new_sdram_controller_grms_wire.addr
		new_sdram_controller_grms_wire_ba    : out   std_logic_vector(1 downto 0);                     --                               .ba
		new_sdram_controller_grms_wire_cas_n : out   std_logic;                                        --                               .cas_n
		new_sdram_controller_grms_wire_cke   : out   std_logic;                                        --                               .cke
		new_sdram_controller_grms_wire_cs_n  : out   std_logic;                                        --                               .cs_n
		new_sdram_controller_grms_wire_dq    : inout std_logic_vector(15 downto 0) := (others => '0'); --                               .dq
		new_sdram_controller_grms_wire_dqm   : out   std_logic_vector(1 downto 0);                     --                               .dqm
		new_sdram_controller_grms_wire_ras_n : out   std_logic;                                        --                               .ras_n
		new_sdram_controller_grms_wire_we_n  : out   std_logic                                         --                               .we_n
	);
end entity p2_grms_qsys;

architecture rtl of p2_grms_qsys is
	component p2_grms_qsys_nios2_qsys_grms is
		port (
			clk                                   : in  std_logic                     := 'X';             -- clk
			reset_n                               : in  std_logic                     := 'X';             -- reset_n
			d_address                             : out std_logic_vector(24 downto 0);                    -- address
			d_byteenable                          : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                                : out std_logic;                                        -- read
			d_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			d_write                               : out std_logic;                                        -- write
			d_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_debug_module_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                             : out std_logic_vector(24 downto 0);                    -- address
			i_read                                : out std_logic;                                        -- read
			i_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			d_irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			jtag_debug_module_resetrequest        : out std_logic;                                        -- reset
			jtag_debug_module_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			jtag_debug_module_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			jtag_debug_module_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			jtag_debug_module_read                : in  std_logic                     := 'X';             -- read
			jtag_debug_module_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			jtag_debug_module_waitrequest         : out std_logic;                                        -- waitrequest
			jtag_debug_module_write               : in  std_logic                     := 'X';             -- write
			jtag_debug_module_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			no_ci_readra                          : out std_logic                                         -- readra
		);
	end component p2_grms_qsys_nios2_qsys_grms;

	component p2_grms_qsys_jtag_uart_grms is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component p2_grms_qsys_jtag_uart_grms;

	component p2_grms_qsys_new_sdram_controller_grms is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(21 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(15 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(11 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(1 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component p2_grms_qsys_new_sdram_controller_grms;

	component p2_grms_qsys_timer_grms is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component p2_grms_qsys_timer_grms;

	component p2_grms_qsys_lcd_16207_grms is
		port (
			reset_n       : in    std_logic                    := 'X';             -- reset_n
			clk           : in    std_logic                    := 'X';             -- clk
			begintransfer : in    std_logic                    := 'X';             -- begintransfer
			read          : in    std_logic                    := 'X';             -- read
			write         : in    std_logic                    := 'X';             -- write
			readdata      : out   std_logic_vector(7 downto 0);                    -- readdata
			writedata     : in    std_logic_vector(7 downto 0) := (others => 'X'); -- writedata
			address       : in    std_logic_vector(1 downto 0) := (others => 'X'); -- address
			LCD_RS        : out   std_logic;                                       -- export
			LCD_RW        : out   std_logic;                                       -- export
			LCD_data      : inout std_logic_vector(7 downto 0) := (others => 'X'); -- export
			LCD_E         : out   std_logic                                        -- export
		);
	end component p2_grms_qsys_lcd_16207_grms;

	component p2_grms_qsys_pa_grms is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(7 downto 0)  := (others => 'X')  -- export
		);
	end component p2_grms_qsys_pa_grms;

	component p2_grms_qsys_pb_grms is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(3 downto 0)  := (others => 'X')  -- export
		);
	end component p2_grms_qsys_pb_grms;

	component p2_grms_qsys_pc_grms is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic                                         -- export
		);
	end component p2_grms_qsys_pc_grms;

	component p2_grms_qsys_pd_grms is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(7 downto 0)                      -- export
		);
	end component p2_grms_qsys_pd_grms;

	component p2_grms_qsys_pf_grms is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(6 downto 0)                      -- export
		);
	end component p2_grms_qsys_pf_grms;

	component p2_grms_qsys_ph_grms is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(3 downto 0)                      -- export
		);
	end component p2_grms_qsys_ph_grms;

	component altera_merlin_master_agent is
		generic (
			PKT_PROTECTION_H          : integer := 80;
			PKT_PROTECTION_L          : integer := 80;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_BURSTWRAP_H           : integer := 79;
			PKT_BURSTWRAP_L           : integer := 77;
			PKT_BURST_SIZE_H          : integer := 86;
			PKT_BURST_SIZE_L          : integer := 84;
			PKT_BURST_TYPE_H          : integer := 94;
			PKT_BURST_TYPE_L          : integer := 93;
			PKT_BYTE_CNT_H            : integer := 76;
			PKT_BYTE_CNT_L            : integer := 74;
			PKT_ADDR_H                : integer := 73;
			PKT_ADDR_L                : integer := 42;
			PKT_TRANS_COMPRESSED_READ : integer := 41;
			PKT_TRANS_POSTED          : integer := 40;
			PKT_TRANS_WRITE           : integer := 39;
			PKT_TRANS_READ            : integer := 38;
			PKT_TRANS_LOCK            : integer := 82;
			PKT_TRANS_EXCLUSIVE       : integer := 83;
			PKT_DATA_H                : integer := 37;
			PKT_DATA_L                : integer := 6;
			PKT_BYTEEN_H              : integer := 5;
			PKT_BYTEEN_L              : integer := 2;
			PKT_SRC_ID_H              : integer := 1;
			PKT_SRC_ID_L              : integer := 1;
			PKT_DEST_ID_H             : integer := 0;
			PKT_DEST_ID_L             : integer := 0;
			PKT_THREAD_ID_H           : integer := 88;
			PKT_THREAD_ID_L           : integer := 87;
			PKT_CACHE_H               : integer := 92;
			PKT_CACHE_L               : integer := 89;
			PKT_DATA_SIDEBAND_H       : integer := 105;
			PKT_DATA_SIDEBAND_L       : integer := 98;
			PKT_QOS_H                 : integer := 109;
			PKT_QOS_L                 : integer := 106;
			PKT_ADDR_SIDEBAND_H       : integer := 97;
			PKT_ADDR_SIDEBAND_L       : integer := 93;
			PKT_RESPONSE_STATUS_H     : integer := 111;
			PKT_RESPONSE_STATUS_L     : integer := 110;
			ST_DATA_W                 : integer := 112;
			ST_CHANNEL_W              : integer := 1;
			AV_BURSTCOUNT_W           : integer := 3;
			SUPPRESS_0_BYTEEN_RSP     : integer := 1;
			ID                        : integer := 1;
			BURSTWRAP_VALUE           : integer := 4;
			CACHE_VALUE               : integer := 0;
			SECURE_ACCESS_BIT         : integer := 1;
			USE_READRESPONSE          : integer := 0;
			USE_WRITERESPONSE         : integer := 0
		);
		port (
			clk                     : in  std_logic                     := 'X';             -- clk
			reset                   : in  std_logic                     := 'X';             -- reset
			av_address              : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			av_write                : in  std_logic                     := 'X';             -- write
			av_read                 : in  std_logic                     := 'X';             -- read
			av_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			av_waitrequest          : out std_logic;                                        -- waitrequest
			av_readdatavalid        : out std_logic;                                        -- readdatavalid
			av_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			av_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			av_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_lock                 : in  std_logic                     := 'X';             -- lock
			cp_valid                : out std_logic;                                        -- valid
			cp_data                 : out std_logic_vector(99 downto 0);                    -- data
			cp_startofpacket        : out std_logic;                                        -- startofpacket
			cp_endofpacket          : out std_logic;                                        -- endofpacket
			cp_ready                : in  std_logic                     := 'X';             -- ready
			rp_valid                : in  std_logic                     := 'X';             -- valid
			rp_data                 : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			rp_channel              : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			rp_startofpacket        : in  std_logic                     := 'X';             -- startofpacket
			rp_endofpacket          : in  std_logic                     := 'X';             -- endofpacket
			rp_ready                : out std_logic;                                        -- ready
			av_response             : out std_logic_vector(1 downto 0);                     -- response
			av_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid   : out std_logic                                         -- writeresponsevalid
		);
	end component altera_merlin_master_agent;

	component p2_grms_qsys_addr_router is
		port (
			sink_ready         : out std_logic;                                        -- ready
			sink_valid         : in  std_logic                     := 'X';             -- valid
			sink_data          : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			src_ready          : in  std_logic                     := 'X';             -- ready
			src_valid          : out std_logic;                                        -- valid
			src_data           : out std_logic_vector(99 downto 0);                    -- data
			src_channel        : out std_logic_vector(13 downto 0);                    -- channel
			src_startofpacket  : out std_logic;                                        -- startofpacket
			src_endofpacket    : out std_logic                                         -- endofpacket
		);
	end component p2_grms_qsys_addr_router;

	component p2_grms_qsys_id_router is
		port (
			sink_ready         : out std_logic;                                        -- ready
			sink_valid         : in  std_logic                     := 'X';             -- valid
			sink_data          : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			src_ready          : in  std_logic                     := 'X';             -- ready
			src_valid          : out std_logic;                                        -- valid
			src_data           : out std_logic_vector(99 downto 0);                    -- data
			src_channel        : out std_logic_vector(13 downto 0);                    -- channel
			src_startofpacket  : out std_logic;                                        -- startofpacket
			src_endofpacket    : out std_logic                                         -- endofpacket
		);
	end component p2_grms_qsys_id_router;

	component p2_grms_qsys_id_router_002 is
		port (
			sink_ready         : out std_logic;                                        -- ready
			sink_valid         : in  std_logic                     := 'X';             -- valid
			sink_data          : in  std_logic_vector(81 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			src_ready          : in  std_logic                     := 'X';             -- ready
			src_valid          : out std_logic;                                        -- valid
			src_data           : out std_logic_vector(81 downto 0);                    -- data
			src_channel        : out std_logic_vector(13 downto 0);                    -- channel
			src_startofpacket  : out std_logic;                                        -- startofpacket
			src_endofpacket    : out std_logic                                         -- endofpacket
		);
	end component p2_grms_qsys_id_router_002;

	component altera_merlin_burst_adapter is
		generic (
			PKT_ADDR_H                : integer := 79;
			PKT_ADDR_L                : integer := 48;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_BYTE_CNT_H            : integer := 5;
			PKT_BYTE_CNT_L            : integer := 0;
			PKT_BYTEEN_H              : integer := 83;
			PKT_BYTEEN_L              : integer := 80;
			PKT_BURST_SIZE_H          : integer := 86;
			PKT_BURST_SIZE_L          : integer := 84;
			PKT_BURST_TYPE_H          : integer := 88;
			PKT_BURST_TYPE_L          : integer := 87;
			PKT_BURSTWRAP_H           : integer := 11;
			PKT_BURSTWRAP_L           : integer := 6;
			PKT_TRANS_COMPRESSED_READ : integer := 14;
			PKT_TRANS_WRITE           : integer := 13;
			PKT_TRANS_READ            : integer := 12;
			OUT_NARROW_SIZE           : integer := 0;
			IN_NARROW_SIZE            : integer := 0;
			OUT_FIXED                 : integer := 0;
			OUT_COMPLETE_WRAP         : integer := 0;
			ST_DATA_W                 : integer := 89;
			ST_CHANNEL_W              : integer := 8;
			OUT_BYTE_CNT_H            : integer := 5;
			OUT_BURSTWRAP_H           : integer := 11;
			COMPRESSED_READ_SUPPORT   : integer := 1;
			BYTEENABLE_SYNTHESIS      : integer := 0;
			PIPE_INPUTS               : integer := 0;
			NO_WRAP_SUPPORT           : integer := 0;
			BURSTWRAP_CONST_MASK      : integer := 0;
			BURSTWRAP_CONST_VALUE     : integer := -1
		);
		port (
			clk                   : in  std_logic                     := 'X';             -- clk
			reset                 : in  std_logic                     := 'X';             -- reset
			sink0_valid           : in  std_logic                     := 'X';             -- valid
			sink0_data            : in  std_logic_vector(81 downto 0) := (others => 'X'); -- data
			sink0_channel         : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			sink0_startofpacket   : in  std_logic                     := 'X';             -- startofpacket
			sink0_endofpacket     : in  std_logic                     := 'X';             -- endofpacket
			sink0_ready           : out std_logic;                                        -- ready
			source0_valid         : out std_logic;                                        -- valid
			source0_data          : out std_logic_vector(81 downto 0);                    -- data
			source0_channel       : out std_logic_vector(13 downto 0);                    -- channel
			source0_startofpacket : out std_logic;                                        -- startofpacket
			source0_endofpacket   : out std_logic;                                        -- endofpacket
			source0_ready         : in  std_logic                     := 'X'              -- ready
		);
	end component altera_merlin_burst_adapter;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS        : integer := 6;
			OUTPUT_RESET_SYNC_EDGES : string  := "deassert";
			SYNC_DEPTH              : integer := 2;
			RESET_REQUEST_PRESENT   : integer := 0
		);
		port (
			reset_in0  : in  std_logic := 'X'; -- reset
			clk        : in  std_logic := 'X'; -- clk
			reset_out  : out std_logic;        -- reset
			reset_req  : out std_logic;        -- reset_req
			reset_in1  : in  std_logic := 'X'; -- reset
			reset_in2  : in  std_logic := 'X'; -- reset
			reset_in3  : in  std_logic := 'X'; -- reset
			reset_in4  : in  std_logic := 'X'; -- reset
			reset_in5  : in  std_logic := 'X'; -- reset
			reset_in6  : in  std_logic := 'X'; -- reset
			reset_in7  : in  std_logic := 'X'; -- reset
			reset_in8  : in  std_logic := 'X'; -- reset
			reset_in9  : in  std_logic := 'X'; -- reset
			reset_in10 : in  std_logic := 'X'; -- reset
			reset_in11 : in  std_logic := 'X'; -- reset
			reset_in12 : in  std_logic := 'X'; -- reset
			reset_in13 : in  std_logic := 'X'; -- reset
			reset_in14 : in  std_logic := 'X'; -- reset
			reset_in15 : in  std_logic := 'X'  -- reset
		);
	end component altera_reset_controller;

	component p2_grms_qsys_cmd_xbar_demux is
		port (
			clk                 : in  std_logic                     := 'X';             -- clk
			reset               : in  std_logic                     := 'X';             -- reset
			sink_ready          : out std_logic;                                        -- ready
			sink_channel        : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			sink_data           : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink_valid          : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- valid
			src0_ready          : in  std_logic                     := 'X';             -- ready
			src0_valid          : out std_logic;                                        -- valid
			src0_data           : out std_logic_vector(99 downto 0);                    -- data
			src0_channel        : out std_logic_vector(13 downto 0);                    -- channel
			src0_startofpacket  : out std_logic;                                        -- startofpacket
			src0_endofpacket    : out std_logic;                                        -- endofpacket
			src1_ready          : in  std_logic                     := 'X';             -- ready
			src1_valid          : out std_logic;                                        -- valid
			src1_data           : out std_logic_vector(99 downto 0);                    -- data
			src1_channel        : out std_logic_vector(13 downto 0);                    -- channel
			src1_startofpacket  : out std_logic;                                        -- startofpacket
			src1_endofpacket    : out std_logic;                                        -- endofpacket
			src2_ready          : in  std_logic                     := 'X';             -- ready
			src2_valid          : out std_logic;                                        -- valid
			src2_data           : out std_logic_vector(99 downto 0);                    -- data
			src2_channel        : out std_logic_vector(13 downto 0);                    -- channel
			src2_startofpacket  : out std_logic;                                        -- startofpacket
			src2_endofpacket    : out std_logic;                                        -- endofpacket
			src3_ready          : in  std_logic                     := 'X';             -- ready
			src3_valid          : out std_logic;                                        -- valid
			src3_data           : out std_logic_vector(99 downto 0);                    -- data
			src3_channel        : out std_logic_vector(13 downto 0);                    -- channel
			src3_startofpacket  : out std_logic;                                        -- startofpacket
			src3_endofpacket    : out std_logic;                                        -- endofpacket
			src4_ready          : in  std_logic                     := 'X';             -- ready
			src4_valid          : out std_logic;                                        -- valid
			src4_data           : out std_logic_vector(99 downto 0);                    -- data
			src4_channel        : out std_logic_vector(13 downto 0);                    -- channel
			src4_startofpacket  : out std_logic;                                        -- startofpacket
			src4_endofpacket    : out std_logic;                                        -- endofpacket
			src5_ready          : in  std_logic                     := 'X';             -- ready
			src5_valid          : out std_logic;                                        -- valid
			src5_data           : out std_logic_vector(99 downto 0);                    -- data
			src5_channel        : out std_logic_vector(13 downto 0);                    -- channel
			src5_startofpacket  : out std_logic;                                        -- startofpacket
			src5_endofpacket    : out std_logic;                                        -- endofpacket
			src6_ready          : in  std_logic                     := 'X';             -- ready
			src6_valid          : out std_logic;                                        -- valid
			src6_data           : out std_logic_vector(99 downto 0);                    -- data
			src6_channel        : out std_logic_vector(13 downto 0);                    -- channel
			src6_startofpacket  : out std_logic;                                        -- startofpacket
			src6_endofpacket    : out std_logic;                                        -- endofpacket
			src7_ready          : in  std_logic                     := 'X';             -- ready
			src7_valid          : out std_logic;                                        -- valid
			src7_data           : out std_logic_vector(99 downto 0);                    -- data
			src7_channel        : out std_logic_vector(13 downto 0);                    -- channel
			src7_startofpacket  : out std_logic;                                        -- startofpacket
			src7_endofpacket    : out std_logic;                                        -- endofpacket
			src8_ready          : in  std_logic                     := 'X';             -- ready
			src8_valid          : out std_logic;                                        -- valid
			src8_data           : out std_logic_vector(99 downto 0);                    -- data
			src8_channel        : out std_logic_vector(13 downto 0);                    -- channel
			src8_startofpacket  : out std_logic;                                        -- startofpacket
			src8_endofpacket    : out std_logic;                                        -- endofpacket
			src9_ready          : in  std_logic                     := 'X';             -- ready
			src9_valid          : out std_logic;                                        -- valid
			src9_data           : out std_logic_vector(99 downto 0);                    -- data
			src9_channel        : out std_logic_vector(13 downto 0);                    -- channel
			src9_startofpacket  : out std_logic;                                        -- startofpacket
			src9_endofpacket    : out std_logic;                                        -- endofpacket
			src10_ready         : in  std_logic                     := 'X';             -- ready
			src10_valid         : out std_logic;                                        -- valid
			src10_data          : out std_logic_vector(99 downto 0);                    -- data
			src10_channel       : out std_logic_vector(13 downto 0);                    -- channel
			src10_startofpacket : out std_logic;                                        -- startofpacket
			src10_endofpacket   : out std_logic;                                        -- endofpacket
			src11_ready         : in  std_logic                     := 'X';             -- ready
			src11_valid         : out std_logic;                                        -- valid
			src11_data          : out std_logic_vector(99 downto 0);                    -- data
			src11_channel       : out std_logic_vector(13 downto 0);                    -- channel
			src11_startofpacket : out std_logic;                                        -- startofpacket
			src11_endofpacket   : out std_logic;                                        -- endofpacket
			src12_ready         : in  std_logic                     := 'X';             -- ready
			src12_valid         : out std_logic;                                        -- valid
			src12_data          : out std_logic_vector(99 downto 0);                    -- data
			src12_channel       : out std_logic_vector(13 downto 0);                    -- channel
			src12_startofpacket : out std_logic;                                        -- startofpacket
			src12_endofpacket   : out std_logic;                                        -- endofpacket
			src13_ready         : in  std_logic                     := 'X';             -- ready
			src13_valid         : out std_logic;                                        -- valid
			src13_data          : out std_logic_vector(99 downto 0);                    -- data
			src13_channel       : out std_logic_vector(13 downto 0);                    -- channel
			src13_startofpacket : out std_logic;                                        -- startofpacket
			src13_endofpacket   : out std_logic                                         -- endofpacket
		);
	end component p2_grms_qsys_cmd_xbar_demux;

	component p2_grms_qsys_cmd_xbar_mux is
		port (
			clk                 : in  std_logic                     := 'X';             -- clk
			reset               : in  std_logic                     := 'X';             -- reset
			src_ready           : in  std_logic                     := 'X';             -- ready
			src_valid           : out std_logic;                                        -- valid
			src_data            : out std_logic_vector(99 downto 0);                    -- data
			src_channel         : out std_logic_vector(13 downto 0);                    -- channel
			src_startofpacket   : out std_logic;                                        -- startofpacket
			src_endofpacket     : out std_logic;                                        -- endofpacket
			sink0_ready         : out std_logic;                                        -- ready
			sink0_valid         : in  std_logic                     := 'X';             -- valid
			sink0_channel       : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			sink0_data          : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink0_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink0_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink1_ready         : out std_logic;                                        -- ready
			sink1_valid         : in  std_logic                     := 'X';             -- valid
			sink1_channel       : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			sink1_data          : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink1_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink1_endofpacket   : in  std_logic                     := 'X'              -- endofpacket
		);
	end component p2_grms_qsys_cmd_xbar_mux;

	component p2_grms_qsys_rsp_xbar_demux is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			sink_ready         : out std_logic;                                        -- ready
			sink_channel       : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- valid
			src0_ready         : in  std_logic                     := 'X';             -- ready
			src0_valid         : out std_logic;                                        -- valid
			src0_data          : out std_logic_vector(99 downto 0);                    -- data
			src0_channel       : out std_logic_vector(13 downto 0);                    -- channel
			src0_startofpacket : out std_logic;                                        -- startofpacket
			src0_endofpacket   : out std_logic;                                        -- endofpacket
			src1_ready         : in  std_logic                     := 'X';             -- ready
			src1_valid         : out std_logic;                                        -- valid
			src1_data          : out std_logic_vector(99 downto 0);                    -- data
			src1_channel       : out std_logic_vector(13 downto 0);                    -- channel
			src1_startofpacket : out std_logic;                                        -- startofpacket
			src1_endofpacket   : out std_logic                                         -- endofpacket
		);
	end component p2_grms_qsys_rsp_xbar_demux;

	component p2_grms_qsys_rsp_xbar_mux is
		port (
			clk                  : in  std_logic                     := 'X';             -- clk
			reset                : in  std_logic                     := 'X';             -- reset
			src_ready            : in  std_logic                     := 'X';             -- ready
			src_valid            : out std_logic;                                        -- valid
			src_data             : out std_logic_vector(99 downto 0);                    -- data
			src_channel          : out std_logic_vector(13 downto 0);                    -- channel
			src_startofpacket    : out std_logic;                                        -- startofpacket
			src_endofpacket      : out std_logic;                                        -- endofpacket
			sink0_ready          : out std_logic;                                        -- ready
			sink0_valid          : in  std_logic                     := 'X';             -- valid
			sink0_channel        : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			sink0_data           : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink0_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink0_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink1_ready          : out std_logic;                                        -- ready
			sink1_valid          : in  std_logic                     := 'X';             -- valid
			sink1_channel        : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			sink1_data           : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink1_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink1_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink2_ready          : out std_logic;                                        -- ready
			sink2_valid          : in  std_logic                     := 'X';             -- valid
			sink2_channel        : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			sink2_data           : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink2_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink2_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink3_ready          : out std_logic;                                        -- ready
			sink3_valid          : in  std_logic                     := 'X';             -- valid
			sink3_channel        : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			sink3_data           : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink3_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink3_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink4_ready          : out std_logic;                                        -- ready
			sink4_valid          : in  std_logic                     := 'X';             -- valid
			sink4_channel        : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			sink4_data           : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink4_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink4_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink5_ready          : out std_logic;                                        -- ready
			sink5_valid          : in  std_logic                     := 'X';             -- valid
			sink5_channel        : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			sink5_data           : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink5_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink5_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink6_ready          : out std_logic;                                        -- ready
			sink6_valid          : in  std_logic                     := 'X';             -- valid
			sink6_channel        : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			sink6_data           : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink6_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink6_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink7_ready          : out std_logic;                                        -- ready
			sink7_valid          : in  std_logic                     := 'X';             -- valid
			sink7_channel        : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			sink7_data           : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink7_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink7_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink8_ready          : out std_logic;                                        -- ready
			sink8_valid          : in  std_logic                     := 'X';             -- valid
			sink8_channel        : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			sink8_data           : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink8_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink8_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink9_ready          : out std_logic;                                        -- ready
			sink9_valid          : in  std_logic                     := 'X';             -- valid
			sink9_channel        : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			sink9_data           : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink9_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink9_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink10_ready         : out std_logic;                                        -- ready
			sink10_valid         : in  std_logic                     := 'X';             -- valid
			sink10_channel       : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			sink10_data          : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink10_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink10_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink11_ready         : out std_logic;                                        -- ready
			sink11_valid         : in  std_logic                     := 'X';             -- valid
			sink11_channel       : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			sink11_data          : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink11_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink11_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink12_ready         : out std_logic;                                        -- ready
			sink12_valid         : in  std_logic                     := 'X';             -- valid
			sink12_channel       : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			sink12_data          : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink12_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink12_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink13_ready         : out std_logic;                                        -- ready
			sink13_valid         : in  std_logic                     := 'X';             -- valid
			sink13_channel       : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			sink13_data          : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink13_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink13_endofpacket   : in  std_logic                     := 'X'              -- endofpacket
		);
	end component p2_grms_qsys_rsp_xbar_mux;

	component p2_grms_qsys_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component p2_grms_qsys_irq_mapper;

	component p2_grms_qsys_nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo is
		generic (
			SYMBOLS_PER_BEAT    : integer := 1;
			BITS_PER_SYMBOL     : integer := 8;
			FIFO_DEPTH          : integer := 16;
			CHANNEL_WIDTH       : integer := 0;
			ERROR_WIDTH         : integer := 0;
			USE_PACKETS         : integer := 0;
			USE_FILL_LEVEL      : integer := 0;
			EMPTY_LATENCY       : integer := 3;
			USE_MEMORY_BLOCKS   : integer := 1;
			USE_STORE_FORWARD   : integer := 0;
			USE_ALMOST_FULL_IF  : integer := 0;
			USE_ALMOST_EMPTY_IF : integer := 0
		);
		port (
			clk               : in  std_logic                      := 'X';             -- clk
			reset             : in  std_logic                      := 'X';             -- reset
			in_data           : in  std_logic_vector(100 downto 0) := (others => 'X'); -- data
			in_valid          : in  std_logic                      := 'X';             -- valid
			in_ready          : out std_logic;                                         -- ready
			in_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			out_data          : out std_logic_vector(100 downto 0);                    -- data
			out_valid         : out std_logic;                                         -- valid
			out_ready         : in  std_logic                      := 'X';             -- ready
			out_startofpacket : out std_logic;                                         -- startofpacket
			out_endofpacket   : out std_logic;                                         -- endofpacket
			csr_address       : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- address
			csr_read          : in  std_logic                      := 'X';             -- read
			csr_write         : in  std_logic                      := 'X';             -- write
			csr_readdata      : out std_logic_vector(31 downto 0);                     -- readdata
			csr_writedata     : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			almost_full_data  : out std_logic;                                         -- data
			almost_empty_data : out std_logic;                                         -- data
			in_empty          : in  std_logic                      := 'X';             -- empty
			out_empty         : out std_logic;                                         -- empty
			in_error          : in  std_logic                      := 'X';             -- error
			out_error         : out std_logic;                                         -- error
			in_channel        : in  std_logic                      := 'X';             -- channel
			out_channel       : out std_logic                                          -- channel
		);
	end component p2_grms_qsys_nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo;

	component p2_grms_qsys_new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo is
		generic (
			SYMBOLS_PER_BEAT    : integer := 1;
			BITS_PER_SYMBOL     : integer := 8;
			FIFO_DEPTH          : integer := 16;
			CHANNEL_WIDTH       : integer := 0;
			ERROR_WIDTH         : integer := 0;
			USE_PACKETS         : integer := 0;
			USE_FILL_LEVEL      : integer := 0;
			EMPTY_LATENCY       : integer := 3;
			USE_MEMORY_BLOCKS   : integer := 1;
			USE_STORE_FORWARD   : integer := 0;
			USE_ALMOST_FULL_IF  : integer := 0;
			USE_ALMOST_EMPTY_IF : integer := 0
		);
		port (
			clk               : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			in_data           : in  std_logic_vector(82 downto 0) := (others => 'X'); -- data
			in_valid          : in  std_logic                     := 'X';             -- valid
			in_ready          : out std_logic;                                        -- ready
			in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			out_data          : out std_logic_vector(82 downto 0);                    -- data
			out_valid         : out std_logic;                                        -- valid
			out_ready         : in  std_logic                     := 'X';             -- ready
			out_startofpacket : out std_logic;                                        -- startofpacket
			out_endofpacket   : out std_logic;                                        -- endofpacket
			csr_address       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			csr_read          : in  std_logic                     := 'X';             -- read
			csr_write         : in  std_logic                     := 'X';             -- write
			csr_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			csr_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			almost_full_data  : out std_logic;                                        -- data
			almost_empty_data : out std_logic;                                        -- data
			in_empty          : in  std_logic                     := 'X';             -- empty
			out_empty         : out std_logic;                                        -- empty
			in_error          : in  std_logic                     := 'X';             -- error
			out_error         : out std_logic;                                        -- error
			in_channel        : in  std_logic                     := 'X';             -- channel
			out_channel       : out std_logic                                         -- channel
		);
	end component p2_grms_qsys_new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo;

	component p2_grms_qsys_new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo is
		generic (
			SYMBOLS_PER_BEAT    : integer := 1;
			BITS_PER_SYMBOL     : integer := 8;
			FIFO_DEPTH          : integer := 16;
			CHANNEL_WIDTH       : integer := 0;
			ERROR_WIDTH         : integer := 0;
			USE_PACKETS         : integer := 0;
			USE_FILL_LEVEL      : integer := 0;
			EMPTY_LATENCY       : integer := 3;
			USE_MEMORY_BLOCKS   : integer := 1;
			USE_STORE_FORWARD   : integer := 0;
			USE_ALMOST_FULL_IF  : integer := 0;
			USE_ALMOST_EMPTY_IF : integer := 0
		);
		port (
			clk               : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			in_data           : in  std_logic_vector(17 downto 0) := (others => 'X'); -- data
			in_valid          : in  std_logic                     := 'X';             -- valid
			in_ready          : out std_logic;                                        -- ready
			out_data          : out std_logic_vector(17 downto 0);                    -- data
			out_valid         : out std_logic;                                        -- valid
			out_ready         : in  std_logic                     := 'X';             -- ready
			csr_address       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			csr_read          : in  std_logic                     := 'X';             -- read
			csr_write         : in  std_logic                     := 'X';             -- write
			csr_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			csr_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			almost_full_data  : out std_logic;                                        -- data
			almost_empty_data : out std_logic;                                        -- data
			in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			out_startofpacket : out std_logic;                                        -- startofpacket
			out_endofpacket   : out std_logic;                                        -- endofpacket
			in_empty          : in  std_logic                     := 'X';             -- empty
			out_empty         : out std_logic;                                        -- empty
			in_error          : in  std_logic                     := 'X';             -- error
			out_error         : out std_logic;                                        -- error
			in_channel        : in  std_logic                     := 'X';             -- channel
			out_channel       : out std_logic                                         -- channel
		);
	end component p2_grms_qsys_new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo;

	component p2_grms_qsys_nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent is
		generic (
			PKT_DATA_H                : integer := 31;
			PKT_DATA_L                : integer := 0;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_SYMBOL_W              : integer := 8;
			PKT_BYTEEN_H              : integer := 71;
			PKT_BYTEEN_L              : integer := 68;
			PKT_ADDR_H                : integer := 63;
			PKT_ADDR_L                : integer := 32;
			PKT_TRANS_COMPRESSED_READ : integer := 67;
			PKT_TRANS_POSTED          : integer := 66;
			PKT_TRANS_WRITE           : integer := 65;
			PKT_TRANS_READ            : integer := 64;
			PKT_TRANS_LOCK            : integer := 87;
			PKT_SRC_ID_H              : integer := 74;
			PKT_SRC_ID_L              : integer := 72;
			PKT_DEST_ID_H             : integer := 77;
			PKT_DEST_ID_L             : integer := 75;
			PKT_BURSTWRAP_H           : integer := 85;
			PKT_BURSTWRAP_L           : integer := 82;
			PKT_BYTE_CNT_H            : integer := 81;
			PKT_BYTE_CNT_L            : integer := 78;
			PKT_PROTECTION_H          : integer := 86;
			PKT_PROTECTION_L          : integer := 86;
			PKT_RESPONSE_STATUS_H     : integer := 89;
			PKT_RESPONSE_STATUS_L     : integer := 88;
			PKT_BURST_SIZE_H          : integer := 92;
			PKT_BURST_SIZE_L          : integer := 90;
			ST_CHANNEL_W              : integer := 8;
			ST_DATA_W                 : integer := 93;
			AVS_BURSTCOUNT_W          : integer := 4;
			SUPPRESS_0_BYTEEN_CMD     : integer := 1;
			PREVENT_FIFO_OVERFLOW     : integer := 0;
			USE_READRESPONSE          : integer := 0;
			USE_WRITERESPONSE         : integer := 0
		);
		port (
			clk                     : in  std_logic                      := 'X';             -- clk
			reset                   : in  std_logic                      := 'X';             -- reset
			m0_address              : out std_logic_vector(24 downto 0);                     -- address
			m0_burstcount           : out std_logic_vector(2 downto 0);                      -- burstcount
			m0_byteenable           : out std_logic_vector(3 downto 0);                      -- byteenable
			m0_debugaccess          : out std_logic;                                         -- debugaccess
			m0_lock                 : out std_logic;                                         -- lock
			m0_readdata             : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                      := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                         -- read
			m0_waitrequest          : in  std_logic                      := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(31 downto 0);                     -- writedata
			m0_write                : out std_logic;                                         -- write
			rp_endofpacket          : out std_logic;                                         -- endofpacket
			rp_ready                : in  std_logic                      := 'X';             -- ready
			rp_valid                : out std_logic;                                         -- valid
			rp_data                 : out std_logic_vector(99 downto 0);                     -- data
			rp_startofpacket        : out std_logic;                                         -- startofpacket
			cp_ready                : out std_logic;                                         -- ready
			cp_valid                : in  std_logic                      := 'X';             -- valid
			cp_data                 : in  std_logic_vector(99 downto 0)  := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                      := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                      := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(13 downto 0)  := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                         -- ready
			rf_sink_valid           : in  std_logic                      := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                      := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                      := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(100 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                      := 'X';             -- ready
			rf_source_valid         : out std_logic;                                         -- valid
			rf_source_startofpacket : out std_logic;                                         -- startofpacket
			rf_source_endofpacket   : out std_logic;                                         -- endofpacket
			rf_source_data          : out std_logic_vector(100 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                         -- ready
			rdata_fifo_sink_valid   : in  std_logic                      := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(33 downto 0)  := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                      := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                         -- valid
			rdata_fifo_src_data     : out std_logic_vector(33 downto 0);                     -- data
			m0_response             : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- response
			m0_writeresponserequest : out std_logic;                                         -- writeresponserequest
			m0_writeresponsevalid   : in  std_logic                      := 'X'              -- writeresponsevalid
		);
	end component p2_grms_qsys_nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent;

	component p2_grms_qsys_new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent is
		generic (
			PKT_DATA_H                : integer := 31;
			PKT_DATA_L                : integer := 0;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_SYMBOL_W              : integer := 8;
			PKT_BYTEEN_H              : integer := 71;
			PKT_BYTEEN_L              : integer := 68;
			PKT_ADDR_H                : integer := 63;
			PKT_ADDR_L                : integer := 32;
			PKT_TRANS_COMPRESSED_READ : integer := 67;
			PKT_TRANS_POSTED          : integer := 66;
			PKT_TRANS_WRITE           : integer := 65;
			PKT_TRANS_READ            : integer := 64;
			PKT_TRANS_LOCK            : integer := 87;
			PKT_SRC_ID_H              : integer := 74;
			PKT_SRC_ID_L              : integer := 72;
			PKT_DEST_ID_H             : integer := 77;
			PKT_DEST_ID_L             : integer := 75;
			PKT_BURSTWRAP_H           : integer := 85;
			PKT_BURSTWRAP_L           : integer := 82;
			PKT_BYTE_CNT_H            : integer := 81;
			PKT_BYTE_CNT_L            : integer := 78;
			PKT_PROTECTION_H          : integer := 86;
			PKT_PROTECTION_L          : integer := 86;
			PKT_RESPONSE_STATUS_H     : integer := 89;
			PKT_RESPONSE_STATUS_L     : integer := 88;
			PKT_BURST_SIZE_H          : integer := 92;
			PKT_BURST_SIZE_L          : integer := 90;
			ST_CHANNEL_W              : integer := 8;
			ST_DATA_W                 : integer := 93;
			AVS_BURSTCOUNT_W          : integer := 4;
			SUPPRESS_0_BYTEEN_CMD     : integer := 1;
			PREVENT_FIFO_OVERFLOW     : integer := 0;
			USE_READRESPONSE          : integer := 0;
			USE_WRITERESPONSE         : integer := 0
		);
		port (
			clk                     : in  std_logic                     := 'X';             -- clk
			reset                   : in  std_logic                     := 'X';             -- reset
			m0_address              : out std_logic_vector(24 downto 0);                    -- address
			m0_burstcount           : out std_logic_vector(1 downto 0);                     -- burstcount
			m0_byteenable           : out std_logic_vector(1 downto 0);                     -- byteenable
			m0_debugaccess          : out std_logic;                                        -- debugaccess
			m0_lock                 : out std_logic;                                        -- lock
			m0_readdata             : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                        -- read
			m0_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(15 downto 0);                    -- writedata
			m0_write                : out std_logic;                                        -- write
			rp_endofpacket          : out std_logic;                                        -- endofpacket
			rp_ready                : in  std_logic                     := 'X';             -- ready
			rp_valid                : out std_logic;                                        -- valid
			rp_data                 : out std_logic_vector(81 downto 0);                    -- data
			rp_startofpacket        : out std_logic;                                        -- startofpacket
			cp_ready                : out std_logic;                                        -- ready
			cp_valid                : in  std_logic                     := 'X';             -- valid
			cp_data                 : in  std_logic_vector(81 downto 0) := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                     := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                     := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                        -- ready
			rf_sink_valid           : in  std_logic                     := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                     := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                     := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(82 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                     := 'X';             -- ready
			rf_source_valid         : out std_logic;                                        -- valid
			rf_source_startofpacket : out std_logic;                                        -- startofpacket
			rf_source_endofpacket   : out std_logic;                                        -- endofpacket
			rf_source_data          : out std_logic_vector(82 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                        -- ready
			rdata_fifo_sink_valid   : in  std_logic                     := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(17 downto 0) := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                     := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                        -- valid
			rdata_fifo_src_data     : out std_logic_vector(17 downto 0);                    -- data
			m0_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			m0_writeresponserequest : out std_logic;                                        -- writeresponserequest
			m0_writeresponsevalid   : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component p2_grms_qsys_new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent;

	component p2_grms_qsys_width_adapter is
		generic (
			IN_PKT_ADDR_H                 : integer := 60;
			IN_PKT_ADDR_L                 : integer := 36;
			IN_PKT_DATA_H                 : integer := 31;
			IN_PKT_DATA_L                 : integer := 0;
			IN_PKT_BYTEEN_H               : integer := 35;
			IN_PKT_BYTEEN_L               : integer := 32;
			IN_PKT_BYTE_CNT_H             : integer := 63;
			IN_PKT_BYTE_CNT_L             : integer := 61;
			IN_PKT_TRANS_COMPRESSED_READ  : integer := 65;
			IN_PKT_BURSTWRAP_H            : integer := 67;
			IN_PKT_BURSTWRAP_L            : integer := 66;
			IN_PKT_BURST_SIZE_H           : integer := 70;
			IN_PKT_BURST_SIZE_L           : integer := 68;
			IN_PKT_RESPONSE_STATUS_H      : integer := 72;
			IN_PKT_RESPONSE_STATUS_L      : integer := 71;
			IN_PKT_TRANS_EXCLUSIVE        : integer := 73;
			IN_PKT_BURST_TYPE_H           : integer := 75;
			IN_PKT_BURST_TYPE_L           : integer := 74;
			IN_ST_DATA_W                  : integer := 76;
			OUT_PKT_ADDR_H                : integer := 60;
			OUT_PKT_ADDR_L                : integer := 36;
			OUT_PKT_DATA_H                : integer := 31;
			OUT_PKT_DATA_L                : integer := 0;
			OUT_PKT_BYTEEN_H              : integer := 35;
			OUT_PKT_BYTEEN_L              : integer := 32;
			OUT_PKT_BYTE_CNT_H            : integer := 63;
			OUT_PKT_BYTE_CNT_L            : integer := 61;
			OUT_PKT_TRANS_COMPRESSED_READ : integer := 65;
			OUT_PKT_BURST_SIZE_H          : integer := 68;
			OUT_PKT_BURST_SIZE_L          : integer := 66;
			OUT_PKT_RESPONSE_STATUS_H     : integer := 70;
			OUT_PKT_RESPONSE_STATUS_L     : integer := 69;
			OUT_PKT_TRANS_EXCLUSIVE       : integer := 71;
			OUT_PKT_BURST_TYPE_H          : integer := 73;
			OUT_PKT_BURST_TYPE_L          : integer := 72;
			OUT_ST_DATA_W                 : integer := 74;
			ST_CHANNEL_W                  : integer := 32;
			OPTIMIZE_FOR_RSP              : integer := 0;
			RESPONSE_PATH                 : integer := 0
		);
		port (
			clk                  : in  std_logic                     := 'X';             -- clk
			reset                : in  std_logic                     := 'X';             -- reset
			in_valid             : in  std_logic                     := 'X';             -- valid
			in_channel           : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			in_startofpacket     : in  std_logic                     := 'X';             -- startofpacket
			in_endofpacket       : in  std_logic                     := 'X';             -- endofpacket
			in_ready             : out std_logic;                                        -- ready
			in_data              : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			out_endofpacket      : out std_logic;                                        -- endofpacket
			out_data             : out std_logic_vector(81 downto 0);                    -- data
			out_channel          : out std_logic_vector(13 downto 0);                    -- channel
			out_valid            : out std_logic;                                        -- valid
			out_ready            : in  std_logic                     := 'X';             -- ready
			out_startofpacket    : out std_logic;                                        -- startofpacket
			in_command_size_data : in  std_logic_vector(2 downto 0)  := (others => 'X')  -- data
		);
	end component p2_grms_qsys_width_adapter;

	component p2_grms_qsys_width_adapter_001 is
		generic (
			IN_PKT_ADDR_H                 : integer := 60;
			IN_PKT_ADDR_L                 : integer := 36;
			IN_PKT_DATA_H                 : integer := 31;
			IN_PKT_DATA_L                 : integer := 0;
			IN_PKT_BYTEEN_H               : integer := 35;
			IN_PKT_BYTEEN_L               : integer := 32;
			IN_PKT_BYTE_CNT_H             : integer := 63;
			IN_PKT_BYTE_CNT_L             : integer := 61;
			IN_PKT_TRANS_COMPRESSED_READ  : integer := 65;
			IN_PKT_BURSTWRAP_H            : integer := 67;
			IN_PKT_BURSTWRAP_L            : integer := 66;
			IN_PKT_BURST_SIZE_H           : integer := 70;
			IN_PKT_BURST_SIZE_L           : integer := 68;
			IN_PKT_RESPONSE_STATUS_H      : integer := 72;
			IN_PKT_RESPONSE_STATUS_L      : integer := 71;
			IN_PKT_TRANS_EXCLUSIVE        : integer := 73;
			IN_PKT_BURST_TYPE_H           : integer := 75;
			IN_PKT_BURST_TYPE_L           : integer := 74;
			IN_ST_DATA_W                  : integer := 76;
			OUT_PKT_ADDR_H                : integer := 60;
			OUT_PKT_ADDR_L                : integer := 36;
			OUT_PKT_DATA_H                : integer := 31;
			OUT_PKT_DATA_L                : integer := 0;
			OUT_PKT_BYTEEN_H              : integer := 35;
			OUT_PKT_BYTEEN_L              : integer := 32;
			OUT_PKT_BYTE_CNT_H            : integer := 63;
			OUT_PKT_BYTE_CNT_L            : integer := 61;
			OUT_PKT_TRANS_COMPRESSED_READ : integer := 65;
			OUT_PKT_BURST_SIZE_H          : integer := 68;
			OUT_PKT_BURST_SIZE_L          : integer := 66;
			OUT_PKT_RESPONSE_STATUS_H     : integer := 70;
			OUT_PKT_RESPONSE_STATUS_L     : integer := 69;
			OUT_PKT_TRANS_EXCLUSIVE       : integer := 71;
			OUT_PKT_BURST_TYPE_H          : integer := 73;
			OUT_PKT_BURST_TYPE_L          : integer := 72;
			OUT_ST_DATA_W                 : integer := 74;
			ST_CHANNEL_W                  : integer := 32;
			OPTIMIZE_FOR_RSP              : integer := 0;
			RESPONSE_PATH                 : integer := 0
		);
		port (
			clk                  : in  std_logic                     := 'X';             -- clk
			reset                : in  std_logic                     := 'X';             -- reset
			in_valid             : in  std_logic                     := 'X';             -- valid
			in_channel           : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			in_startofpacket     : in  std_logic                     := 'X';             -- startofpacket
			in_endofpacket       : in  std_logic                     := 'X';             -- endofpacket
			in_ready             : out std_logic;                                        -- ready
			in_data              : in  std_logic_vector(81 downto 0) := (others => 'X'); -- data
			out_endofpacket      : out std_logic;                                        -- endofpacket
			out_data             : out std_logic_vector(99 downto 0);                    -- data
			out_channel          : out std_logic_vector(13 downto 0);                    -- channel
			out_valid            : out std_logic;                                        -- valid
			out_ready            : in  std_logic                     := 'X';             -- ready
			out_startofpacket    : out std_logic;                                        -- startofpacket
			in_command_size_data : in  std_logic_vector(2 downto 0)  := (others => 'X')  -- data
		);
	end component p2_grms_qsys_width_adapter_001;

	component p2_grms_qsys_nios2_qsys_grms_instruction_master_translator is
		generic (
			AV_ADDRESS_W                : integer := 32;
			AV_DATA_W                   : integer := 32;
			AV_BURSTCOUNT_W             : integer := 4;
			AV_BYTEENABLE_W             : integer := 4;
			UAV_ADDRESS_W               : integer := 38;
			UAV_BURSTCOUNT_W            : integer := 10;
			USE_READ                    : integer := 1;
			USE_WRITE                   : integer := 1;
			USE_BEGINBURSTTRANSFER      : integer := 0;
			USE_BEGINTRANSFER           : integer := 0;
			USE_CHIPSELECT              : integer := 0;
			USE_BURSTCOUNT              : integer := 1;
			USE_READDATAVALID           : integer := 1;
			USE_WAITREQUEST             : integer := 1;
			USE_READRESPONSE            : integer := 0;
			USE_WRITERESPONSE           : integer := 0;
			AV_SYMBOLS_PER_WORD         : integer := 4;
			AV_ADDRESS_SYMBOLS          : integer := 0;
			AV_BURSTCOUNT_SYMBOLS       : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR  : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR : integer := 0;
			AV_LINEWRAPBURSTS           : integer := 0;
			AV_REGISTERINCOMINGSIGNALS  : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : out std_logic_vector(24 downto 0);                    -- address
			uav_burstcount           : out std_logic_vector(2 downto 0);                     -- burstcount
			uav_read                 : out std_logic;                                        -- read
			uav_write                : out std_logic;                                        -- write
			uav_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			uav_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			uav_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			uav_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			uav_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			uav_lock                 : out std_logic;                                        -- lock
			uav_debugaccess          : out std_logic;                                        -- debugaccess
			av_address               : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			av_waitrequest           : out std_logic;                                        -- waitrequest
			av_read                  : in  std_logic                     := 'X';             -- read
			av_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			av_burstcount            : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			av_byteenable            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			av_beginbursttransfer    : in  std_logic                     := 'X';             -- beginbursttransfer
			av_begintransfer         : in  std_logic                     := 'X';             -- begintransfer
			av_chipselect            : in  std_logic                     := 'X';             -- chipselect
			av_readdatavalid         : out std_logic;                                        -- readdatavalid
			av_write                 : in  std_logic                     := 'X';             -- write
			av_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_lock                  : in  std_logic                     := 'X';             -- lock
			av_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			uav_clken                : out std_logic;                                        -- clken
			av_clken                 : in  std_logic                     := 'X';             -- clken
			uav_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			av_response              : out std_logic_vector(1 downto 0);                     -- response
			uav_writeresponserequest : out std_logic;                                        -- writeresponserequest
			uav_writeresponsevalid   : in  std_logic                     := 'X';             -- writeresponsevalid
			av_writeresponserequest  : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid    : out std_logic                                         -- writeresponsevalid
		);
	end component p2_grms_qsys_nios2_qsys_grms_instruction_master_translator;

	component p2_grms_qsys_nios2_qsys_grms_data_master_translator is
		generic (
			AV_ADDRESS_W                : integer := 32;
			AV_DATA_W                   : integer := 32;
			AV_BURSTCOUNT_W             : integer := 4;
			AV_BYTEENABLE_W             : integer := 4;
			UAV_ADDRESS_W               : integer := 38;
			UAV_BURSTCOUNT_W            : integer := 10;
			USE_READ                    : integer := 1;
			USE_WRITE                   : integer := 1;
			USE_BEGINBURSTTRANSFER      : integer := 0;
			USE_BEGINTRANSFER           : integer := 0;
			USE_CHIPSELECT              : integer := 0;
			USE_BURSTCOUNT              : integer := 1;
			USE_READDATAVALID           : integer := 1;
			USE_WAITREQUEST             : integer := 1;
			USE_READRESPONSE            : integer := 0;
			USE_WRITERESPONSE           : integer := 0;
			AV_SYMBOLS_PER_WORD         : integer := 4;
			AV_ADDRESS_SYMBOLS          : integer := 0;
			AV_BURSTCOUNT_SYMBOLS       : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR  : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR : integer := 0;
			AV_LINEWRAPBURSTS           : integer := 0;
			AV_REGISTERINCOMINGSIGNALS  : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : out std_logic_vector(24 downto 0);                    -- address
			uav_burstcount           : out std_logic_vector(2 downto 0);                     -- burstcount
			uav_read                 : out std_logic;                                        -- read
			uav_write                : out std_logic;                                        -- write
			uav_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			uav_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			uav_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			uav_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			uav_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			uav_lock                 : out std_logic;                                        -- lock
			uav_debugaccess          : out std_logic;                                        -- debugaccess
			av_address               : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			av_waitrequest           : out std_logic;                                        -- waitrequest
			av_byteenable            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			av_read                  : in  std_logic                     := 'X';             -- read
			av_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			av_write                 : in  std_logic                     := 'X';             -- write
			av_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			av_burstcount            : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			av_beginbursttransfer    : in  std_logic                     := 'X';             -- beginbursttransfer
			av_begintransfer         : in  std_logic                     := 'X';             -- begintransfer
			av_chipselect            : in  std_logic                     := 'X';             -- chipselect
			av_readdatavalid         : out std_logic;                                        -- readdatavalid
			av_lock                  : in  std_logic                     := 'X';             -- lock
			uav_clken                : out std_logic;                                        -- clken
			av_clken                 : in  std_logic                     := 'X';             -- clken
			uav_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			av_response              : out std_logic_vector(1 downto 0);                     -- response
			uav_writeresponserequest : out std_logic;                                        -- writeresponserequest
			uav_writeresponsevalid   : in  std_logic                     := 'X';             -- writeresponsevalid
			av_writeresponserequest  : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid    : out std_logic                                         -- writeresponsevalid
		);
	end component p2_grms_qsys_nios2_qsys_grms_data_master_translator;

	component p2_grms_qsys_nios2_qsys_grms_jtag_debug_module_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(8 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_writebyteenable       : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component p2_grms_qsys_nios2_qsys_grms_jtag_debug_module_translator;

	component p2_grms_qsys_jtag_uart_grms_avalon_jtag_slave_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(0 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_chipselect            : out std_logic;                                        -- chipselect
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_writebyteenable       : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component p2_grms_qsys_jtag_uart_grms_avalon_jtag_slave_translator;

	component p2_grms_qsys_new_sdram_controller_grms_s1_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(15 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(21 downto 0);                    -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(15 downto 0);                    -- writedata
			av_byteenable            : out std_logic_vector(1 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_chipselect            : out std_logic;                                        -- chipselect
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_writebyteenable       : out std_logic_vector(1 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component p2_grms_qsys_new_sdram_controller_grms_s1_translator;

	component p2_grms_qsys_timer_grms_s1_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(2 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_readdata              : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(15 downto 0);                    -- writedata
			av_chipselect            : out std_logic;                                        -- chipselect
			av_read                  : out std_logic;                                        -- read
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component p2_grms_qsys_timer_grms_s1_translator;

	component p2_grms_qsys_lcd_16207_grms_control_slave_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(1 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(7 downto 0);                     -- writedata
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component p2_grms_qsys_lcd_16207_grms_control_slave_translator;

	component p2_grms_qsys_pa_grms_s1_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(1 downto 0);                     -- address
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component p2_grms_qsys_pa_grms_s1_translator;

	component p2_grms_qsys_pc_grms_s1_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(1 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_chipselect            : out std_logic;                                        -- chipselect
			av_read                  : out std_logic;                                        -- read
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component p2_grms_qsys_pc_grms_s1_translator;

	signal nios2_qsys_grms_instruction_master_waitrequest                                                         : std_logic;                      -- nios2_qsys_grms_instruction_master_translator:av_waitrequest -> nios2_qsys_grms:i_waitrequest
	signal nios2_qsys_grms_instruction_master_address                                                             : std_logic_vector(24 downto 0);  -- nios2_qsys_grms:i_address -> nios2_qsys_grms_instruction_master_translator:av_address
	signal nios2_qsys_grms_instruction_master_read                                                                : std_logic;                      -- nios2_qsys_grms:i_read -> nios2_qsys_grms_instruction_master_translator:av_read
	signal nios2_qsys_grms_instruction_master_readdata                                                            : std_logic_vector(31 downto 0);  -- nios2_qsys_grms_instruction_master_translator:av_readdata -> nios2_qsys_grms:i_readdata
	signal nios2_qsys_grms_data_master_waitrequest                                                                : std_logic;                      -- nios2_qsys_grms_data_master_translator:av_waitrequest -> nios2_qsys_grms:d_waitrequest
	signal nios2_qsys_grms_data_master_writedata                                                                  : std_logic_vector(31 downto 0);  -- nios2_qsys_grms:d_writedata -> nios2_qsys_grms_data_master_translator:av_writedata
	signal nios2_qsys_grms_data_master_address                                                                    : std_logic_vector(24 downto 0);  -- nios2_qsys_grms:d_address -> nios2_qsys_grms_data_master_translator:av_address
	signal nios2_qsys_grms_data_master_write                                                                      : std_logic;                      -- nios2_qsys_grms:d_write -> nios2_qsys_grms_data_master_translator:av_write
	signal nios2_qsys_grms_data_master_read                                                                       : std_logic;                      -- nios2_qsys_grms:d_read -> nios2_qsys_grms_data_master_translator:av_read
	signal nios2_qsys_grms_data_master_readdata                                                                   : std_logic_vector(31 downto 0);  -- nios2_qsys_grms_data_master_translator:av_readdata -> nios2_qsys_grms:d_readdata
	signal nios2_qsys_grms_data_master_debugaccess                                                                : std_logic;                      -- nios2_qsys_grms:jtag_debug_module_debugaccess_to_roms -> nios2_qsys_grms_data_master_translator:av_debugaccess
	signal nios2_qsys_grms_data_master_byteenable                                                                 : std_logic_vector(3 downto 0);   -- nios2_qsys_grms:d_byteenable -> nios2_qsys_grms_data_master_translator:av_byteenable
	signal nios2_qsys_grms_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest                           : std_logic;                      -- nios2_qsys_grms:jtag_debug_module_waitrequest -> nios2_qsys_grms_jtag_debug_module_translator:av_waitrequest
	signal nios2_qsys_grms_jtag_debug_module_translator_avalon_anti_slave_0_writedata                             : std_logic_vector(31 downto 0);  -- nios2_qsys_grms_jtag_debug_module_translator:av_writedata -> nios2_qsys_grms:jtag_debug_module_writedata
	signal nios2_qsys_grms_jtag_debug_module_translator_avalon_anti_slave_0_address                               : std_logic_vector(8 downto 0);   -- nios2_qsys_grms_jtag_debug_module_translator:av_address -> nios2_qsys_grms:jtag_debug_module_address
	signal nios2_qsys_grms_jtag_debug_module_translator_avalon_anti_slave_0_write                                 : std_logic;                      -- nios2_qsys_grms_jtag_debug_module_translator:av_write -> nios2_qsys_grms:jtag_debug_module_write
	signal nios2_qsys_grms_jtag_debug_module_translator_avalon_anti_slave_0_read                                  : std_logic;                      -- nios2_qsys_grms_jtag_debug_module_translator:av_read -> nios2_qsys_grms:jtag_debug_module_read
	signal nios2_qsys_grms_jtag_debug_module_translator_avalon_anti_slave_0_readdata                              : std_logic_vector(31 downto 0);  -- nios2_qsys_grms:jtag_debug_module_readdata -> nios2_qsys_grms_jtag_debug_module_translator:av_readdata
	signal nios2_qsys_grms_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess                           : std_logic;                      -- nios2_qsys_grms_jtag_debug_module_translator:av_debugaccess -> nios2_qsys_grms:jtag_debug_module_debugaccess
	signal nios2_qsys_grms_jtag_debug_module_translator_avalon_anti_slave_0_byteenable                            : std_logic_vector(3 downto 0);   -- nios2_qsys_grms_jtag_debug_module_translator:av_byteenable -> nios2_qsys_grms:jtag_debug_module_byteenable
	signal jtag_uart_grms_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest                            : std_logic;                      -- jtag_uart_grms:av_waitrequest -> jtag_uart_grms_avalon_jtag_slave_translator:av_waitrequest
	signal jtag_uart_grms_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata                              : std_logic_vector(31 downto 0);  -- jtag_uart_grms_avalon_jtag_slave_translator:av_writedata -> jtag_uart_grms:av_writedata
	signal jtag_uart_grms_avalon_jtag_slave_translator_avalon_anti_slave_0_address                                : std_logic_vector(0 downto 0);   -- jtag_uart_grms_avalon_jtag_slave_translator:av_address -> jtag_uart_grms:av_address
	signal jtag_uart_grms_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect                             : std_logic;                      -- jtag_uart_grms_avalon_jtag_slave_translator:av_chipselect -> jtag_uart_grms:av_chipselect
	signal jtag_uart_grms_avalon_jtag_slave_translator_avalon_anti_slave_0_write                                  : std_logic;                      -- jtag_uart_grms_avalon_jtag_slave_translator:av_write -> jtag_uart_grms_avalon_jtag_slave_translator_avalon_anti_slave_0_write:in
	signal jtag_uart_grms_avalon_jtag_slave_translator_avalon_anti_slave_0_read                                   : std_logic;                      -- jtag_uart_grms_avalon_jtag_slave_translator:av_read -> jtag_uart_grms_avalon_jtag_slave_translator_avalon_anti_slave_0_read:in
	signal jtag_uart_grms_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata                               : std_logic_vector(31 downto 0);  -- jtag_uart_grms:av_readdata -> jtag_uart_grms_avalon_jtag_slave_translator:av_readdata
	signal new_sdram_controller_grms_s1_translator_avalon_anti_slave_0_waitrequest                                : std_logic;                      -- new_sdram_controller_grms:za_waitrequest -> new_sdram_controller_grms_s1_translator:av_waitrequest
	signal new_sdram_controller_grms_s1_translator_avalon_anti_slave_0_writedata                                  : std_logic_vector(15 downto 0);  -- new_sdram_controller_grms_s1_translator:av_writedata -> new_sdram_controller_grms:az_data
	signal new_sdram_controller_grms_s1_translator_avalon_anti_slave_0_address                                    : std_logic_vector(21 downto 0);  -- new_sdram_controller_grms_s1_translator:av_address -> new_sdram_controller_grms:az_addr
	signal new_sdram_controller_grms_s1_translator_avalon_anti_slave_0_chipselect                                 : std_logic;                      -- new_sdram_controller_grms_s1_translator:av_chipselect -> new_sdram_controller_grms:az_cs
	signal new_sdram_controller_grms_s1_translator_avalon_anti_slave_0_write                                      : std_logic;                      -- new_sdram_controller_grms_s1_translator:av_write -> new_sdram_controller_grms_s1_translator_avalon_anti_slave_0_write:in
	signal new_sdram_controller_grms_s1_translator_avalon_anti_slave_0_read                                       : std_logic;                      -- new_sdram_controller_grms_s1_translator:av_read -> new_sdram_controller_grms_s1_translator_avalon_anti_slave_0_read:in
	signal new_sdram_controller_grms_s1_translator_avalon_anti_slave_0_readdata                                   : std_logic_vector(15 downto 0);  -- new_sdram_controller_grms:za_data -> new_sdram_controller_grms_s1_translator:av_readdata
	signal new_sdram_controller_grms_s1_translator_avalon_anti_slave_0_readdatavalid                              : std_logic;                      -- new_sdram_controller_grms:za_valid -> new_sdram_controller_grms_s1_translator:av_readdatavalid
	signal new_sdram_controller_grms_s1_translator_avalon_anti_slave_0_byteenable                                 : std_logic_vector(1 downto 0);   -- new_sdram_controller_grms_s1_translator:av_byteenable -> new_sdram_controller_grms_s1_translator_avalon_anti_slave_0_byteenable:in
	signal timer_grms_s1_translator_avalon_anti_slave_0_writedata                                                 : std_logic_vector(15 downto 0);  -- timer_grms_s1_translator:av_writedata -> timer_grms:writedata
	signal timer_grms_s1_translator_avalon_anti_slave_0_address                                                   : std_logic_vector(2 downto 0);   -- timer_grms_s1_translator:av_address -> timer_grms:address
	signal timer_grms_s1_translator_avalon_anti_slave_0_chipselect                                                : std_logic;                      -- timer_grms_s1_translator:av_chipselect -> timer_grms:chipselect
	signal timer_grms_s1_translator_avalon_anti_slave_0_write                                                     : std_logic;                      -- timer_grms_s1_translator:av_write -> timer_grms_s1_translator_avalon_anti_slave_0_write:in
	signal timer_grms_s1_translator_avalon_anti_slave_0_readdata                                                  : std_logic_vector(15 downto 0);  -- timer_grms:readdata -> timer_grms_s1_translator:av_readdata
	signal lcd_16207_grms_control_slave_translator_avalon_anti_slave_0_writedata                                  : std_logic_vector(7 downto 0);   -- lcd_16207_grms_control_slave_translator:av_writedata -> lcd_16207_grms:writedata
	signal lcd_16207_grms_control_slave_translator_avalon_anti_slave_0_address                                    : std_logic_vector(1 downto 0);   -- lcd_16207_grms_control_slave_translator:av_address -> lcd_16207_grms:address
	signal lcd_16207_grms_control_slave_translator_avalon_anti_slave_0_write                                      : std_logic;                      -- lcd_16207_grms_control_slave_translator:av_write -> lcd_16207_grms:write
	signal lcd_16207_grms_control_slave_translator_avalon_anti_slave_0_read                                       : std_logic;                      -- lcd_16207_grms_control_slave_translator:av_read -> lcd_16207_grms:read
	signal lcd_16207_grms_control_slave_translator_avalon_anti_slave_0_readdata                                   : std_logic_vector(7 downto 0);   -- lcd_16207_grms:readdata -> lcd_16207_grms_control_slave_translator:av_readdata
	signal lcd_16207_grms_control_slave_translator_avalon_anti_slave_0_begintransfer                              : std_logic;                      -- lcd_16207_grms_control_slave_translator:av_begintransfer -> lcd_16207_grms:begintransfer
	signal pa_grms_s1_translator_avalon_anti_slave_0_address                                                      : std_logic_vector(1 downto 0);   -- pa_grms_s1_translator:av_address -> pa_grms:address
	signal pa_grms_s1_translator_avalon_anti_slave_0_readdata                                                     : std_logic_vector(31 downto 0);  -- pa_grms:readdata -> pa_grms_s1_translator:av_readdata
	signal pb_grms_s1_translator_avalon_anti_slave_0_address                                                      : std_logic_vector(1 downto 0);   -- pb_grms_s1_translator:av_address -> pb_grms:address
	signal pb_grms_s1_translator_avalon_anti_slave_0_readdata                                                     : std_logic_vector(31 downto 0);  -- pb_grms:readdata -> pb_grms_s1_translator:av_readdata
	signal pc_grms_s1_translator_avalon_anti_slave_0_writedata                                                    : std_logic_vector(31 downto 0);  -- pc_grms_s1_translator:av_writedata -> pc_grms:writedata
	signal pc_grms_s1_translator_avalon_anti_slave_0_address                                                      : std_logic_vector(1 downto 0);   -- pc_grms_s1_translator:av_address -> pc_grms:address
	signal pc_grms_s1_translator_avalon_anti_slave_0_chipselect                                                   : std_logic;                      -- pc_grms_s1_translator:av_chipselect -> pc_grms:chipselect
	signal pc_grms_s1_translator_avalon_anti_slave_0_write                                                        : std_logic;                      -- pc_grms_s1_translator:av_write -> pc_grms_s1_translator_avalon_anti_slave_0_write:in
	signal pc_grms_s1_translator_avalon_anti_slave_0_readdata                                                     : std_logic_vector(31 downto 0);  -- pc_grms:readdata -> pc_grms_s1_translator:av_readdata
	signal pd_grms_s1_translator_avalon_anti_slave_0_writedata                                                    : std_logic_vector(31 downto 0);  -- pd_grms_s1_translator:av_writedata -> pd_grms:writedata
	signal pd_grms_s1_translator_avalon_anti_slave_0_address                                                      : std_logic_vector(1 downto 0);   -- pd_grms_s1_translator:av_address -> pd_grms:address
	signal pd_grms_s1_translator_avalon_anti_slave_0_chipselect                                                   : std_logic;                      -- pd_grms_s1_translator:av_chipselect -> pd_grms:chipselect
	signal pd_grms_s1_translator_avalon_anti_slave_0_write                                                        : std_logic;                      -- pd_grms_s1_translator:av_write -> pd_grms_s1_translator_avalon_anti_slave_0_write:in
	signal pd_grms_s1_translator_avalon_anti_slave_0_readdata                                                     : std_logic_vector(31 downto 0);  -- pd_grms:readdata -> pd_grms_s1_translator:av_readdata
	signal pe_grms_s1_translator_avalon_anti_slave_0_writedata                                                    : std_logic_vector(31 downto 0);  -- pe_grms_s1_translator:av_writedata -> pe_grms:writedata
	signal pe_grms_s1_translator_avalon_anti_slave_0_address                                                      : std_logic_vector(1 downto 0);   -- pe_grms_s1_translator:av_address -> pe_grms:address
	signal pe_grms_s1_translator_avalon_anti_slave_0_chipselect                                                   : std_logic;                      -- pe_grms_s1_translator:av_chipselect -> pe_grms:chipselect
	signal pe_grms_s1_translator_avalon_anti_slave_0_write                                                        : std_logic;                      -- pe_grms_s1_translator:av_write -> pe_grms_s1_translator_avalon_anti_slave_0_write:in
	signal pe_grms_s1_translator_avalon_anti_slave_0_readdata                                                     : std_logic_vector(31 downto 0);  -- pe_grms:readdata -> pe_grms_s1_translator:av_readdata
	signal pf_grms_s1_translator_avalon_anti_slave_0_writedata                                                    : std_logic_vector(31 downto 0);  -- pf_grms_s1_translator:av_writedata -> pf_grms:writedata
	signal pf_grms_s1_translator_avalon_anti_slave_0_address                                                      : std_logic_vector(1 downto 0);   -- pf_grms_s1_translator:av_address -> pf_grms:address
	signal pf_grms_s1_translator_avalon_anti_slave_0_chipselect                                                   : std_logic;                      -- pf_grms_s1_translator:av_chipselect -> pf_grms:chipselect
	signal pf_grms_s1_translator_avalon_anti_slave_0_write                                                        : std_logic;                      -- pf_grms_s1_translator:av_write -> pf_grms_s1_translator_avalon_anti_slave_0_write:in
	signal pf_grms_s1_translator_avalon_anti_slave_0_readdata                                                     : std_logic_vector(31 downto 0);  -- pf_grms:readdata -> pf_grms_s1_translator:av_readdata
	signal pg_grms_s1_translator_avalon_anti_slave_0_writedata                                                    : std_logic_vector(31 downto 0);  -- pg_grms_s1_translator:av_writedata -> pg_grms:writedata
	signal pg_grms_s1_translator_avalon_anti_slave_0_address                                                      : std_logic_vector(1 downto 0);   -- pg_grms_s1_translator:av_address -> pg_grms:address
	signal pg_grms_s1_translator_avalon_anti_slave_0_chipselect                                                   : std_logic;                      -- pg_grms_s1_translator:av_chipselect -> pg_grms:chipselect
	signal pg_grms_s1_translator_avalon_anti_slave_0_write                                                        : std_logic;                      -- pg_grms_s1_translator:av_write -> pg_grms_s1_translator_avalon_anti_slave_0_write:in
	signal pg_grms_s1_translator_avalon_anti_slave_0_readdata                                                     : std_logic_vector(31 downto 0);  -- pg_grms:readdata -> pg_grms_s1_translator:av_readdata
	signal ph_grms_s1_translator_avalon_anti_slave_0_writedata                                                    : std_logic_vector(31 downto 0);  -- ph_grms_s1_translator:av_writedata -> ph_grms:writedata
	signal ph_grms_s1_translator_avalon_anti_slave_0_address                                                      : std_logic_vector(1 downto 0);   -- ph_grms_s1_translator:av_address -> ph_grms:address
	signal ph_grms_s1_translator_avalon_anti_slave_0_chipselect                                                   : std_logic;                      -- ph_grms_s1_translator:av_chipselect -> ph_grms:chipselect
	signal ph_grms_s1_translator_avalon_anti_slave_0_write                                                        : std_logic;                      -- ph_grms_s1_translator:av_write -> ph_grms_s1_translator_avalon_anti_slave_0_write:in
	signal ph_grms_s1_translator_avalon_anti_slave_0_readdata                                                     : std_logic_vector(31 downto 0);  -- ph_grms:readdata -> ph_grms_s1_translator:av_readdata
	signal pi_grms_s1_translator_avalon_anti_slave_0_writedata                                                    : std_logic_vector(31 downto 0);  -- pi_grms_s1_translator:av_writedata -> pi_grms:writedata
	signal pi_grms_s1_translator_avalon_anti_slave_0_address                                                      : std_logic_vector(1 downto 0);   -- pi_grms_s1_translator:av_address -> pi_grms:address
	signal pi_grms_s1_translator_avalon_anti_slave_0_chipselect                                                   : std_logic;                      -- pi_grms_s1_translator:av_chipselect -> pi_grms:chipselect
	signal pi_grms_s1_translator_avalon_anti_slave_0_write                                                        : std_logic;                      -- pi_grms_s1_translator:av_write -> pi_grms_s1_translator_avalon_anti_slave_0_write:in
	signal pi_grms_s1_translator_avalon_anti_slave_0_readdata                                                     : std_logic_vector(31 downto 0);  -- pi_grms:readdata -> pi_grms_s1_translator:av_readdata
	signal nios2_qsys_grms_instruction_master_translator_avalon_universal_master_0_waitrequest                    : std_logic;                      -- nios2_qsys_grms_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios2_qsys_grms_instruction_master_translator:uav_waitrequest
	signal nios2_qsys_grms_instruction_master_translator_avalon_universal_master_0_burstcount                     : std_logic_vector(2 downto 0);   -- nios2_qsys_grms_instruction_master_translator:uav_burstcount -> nios2_qsys_grms_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	signal nios2_qsys_grms_instruction_master_translator_avalon_universal_master_0_writedata                      : std_logic_vector(31 downto 0);  -- nios2_qsys_grms_instruction_master_translator:uav_writedata -> nios2_qsys_grms_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	signal nios2_qsys_grms_instruction_master_translator_avalon_universal_master_0_address                        : std_logic_vector(24 downto 0);  -- nios2_qsys_grms_instruction_master_translator:uav_address -> nios2_qsys_grms_instruction_master_translator_avalon_universal_master_0_agent:av_address
	signal nios2_qsys_grms_instruction_master_translator_avalon_universal_master_0_lock                           : std_logic;                      -- nios2_qsys_grms_instruction_master_translator:uav_lock -> nios2_qsys_grms_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	signal nios2_qsys_grms_instruction_master_translator_avalon_universal_master_0_write                          : std_logic;                      -- nios2_qsys_grms_instruction_master_translator:uav_write -> nios2_qsys_grms_instruction_master_translator_avalon_universal_master_0_agent:av_write
	signal nios2_qsys_grms_instruction_master_translator_avalon_universal_master_0_read                           : std_logic;                      -- nios2_qsys_grms_instruction_master_translator:uav_read -> nios2_qsys_grms_instruction_master_translator_avalon_universal_master_0_agent:av_read
	signal nios2_qsys_grms_instruction_master_translator_avalon_universal_master_0_readdata                       : std_logic_vector(31 downto 0);  -- nios2_qsys_grms_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> nios2_qsys_grms_instruction_master_translator:uav_readdata
	signal nios2_qsys_grms_instruction_master_translator_avalon_universal_master_0_debugaccess                    : std_logic;                      -- nios2_qsys_grms_instruction_master_translator:uav_debugaccess -> nios2_qsys_grms_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	signal nios2_qsys_grms_instruction_master_translator_avalon_universal_master_0_byteenable                     : std_logic_vector(3 downto 0);   -- nios2_qsys_grms_instruction_master_translator:uav_byteenable -> nios2_qsys_grms_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	signal nios2_qsys_grms_instruction_master_translator_avalon_universal_master_0_readdatavalid                  : std_logic;                      -- nios2_qsys_grms_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios2_qsys_grms_instruction_master_translator:uav_readdatavalid
	signal nios2_qsys_grms_data_master_translator_avalon_universal_master_0_waitrequest                           : std_logic;                      -- nios2_qsys_grms_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios2_qsys_grms_data_master_translator:uav_waitrequest
	signal nios2_qsys_grms_data_master_translator_avalon_universal_master_0_burstcount                            : std_logic_vector(2 downto 0);   -- nios2_qsys_grms_data_master_translator:uav_burstcount -> nios2_qsys_grms_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	signal nios2_qsys_grms_data_master_translator_avalon_universal_master_0_writedata                             : std_logic_vector(31 downto 0);  -- nios2_qsys_grms_data_master_translator:uav_writedata -> nios2_qsys_grms_data_master_translator_avalon_universal_master_0_agent:av_writedata
	signal nios2_qsys_grms_data_master_translator_avalon_universal_master_0_address                               : std_logic_vector(24 downto 0);  -- nios2_qsys_grms_data_master_translator:uav_address -> nios2_qsys_grms_data_master_translator_avalon_universal_master_0_agent:av_address
	signal nios2_qsys_grms_data_master_translator_avalon_universal_master_0_lock                                  : std_logic;                      -- nios2_qsys_grms_data_master_translator:uav_lock -> nios2_qsys_grms_data_master_translator_avalon_universal_master_0_agent:av_lock
	signal nios2_qsys_grms_data_master_translator_avalon_universal_master_0_write                                 : std_logic;                      -- nios2_qsys_grms_data_master_translator:uav_write -> nios2_qsys_grms_data_master_translator_avalon_universal_master_0_agent:av_write
	signal nios2_qsys_grms_data_master_translator_avalon_universal_master_0_read                                  : std_logic;                      -- nios2_qsys_grms_data_master_translator:uav_read -> nios2_qsys_grms_data_master_translator_avalon_universal_master_0_agent:av_read
	signal nios2_qsys_grms_data_master_translator_avalon_universal_master_0_readdata                              : std_logic_vector(31 downto 0);  -- nios2_qsys_grms_data_master_translator_avalon_universal_master_0_agent:av_readdata -> nios2_qsys_grms_data_master_translator:uav_readdata
	signal nios2_qsys_grms_data_master_translator_avalon_universal_master_0_debugaccess                           : std_logic;                      -- nios2_qsys_grms_data_master_translator:uav_debugaccess -> nios2_qsys_grms_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	signal nios2_qsys_grms_data_master_translator_avalon_universal_master_0_byteenable                            : std_logic_vector(3 downto 0);   -- nios2_qsys_grms_data_master_translator:uav_byteenable -> nios2_qsys_grms_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	signal nios2_qsys_grms_data_master_translator_avalon_universal_master_0_readdatavalid                         : std_logic;                      -- nios2_qsys_grms_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios2_qsys_grms_data_master_translator:uav_readdatavalid
	signal nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest             : std_logic;                      -- nios2_qsys_grms_jtag_debug_module_translator:uav_waitrequest -> nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount              : std_logic_vector(2 downto 0);   -- nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> nios2_qsys_grms_jtag_debug_module_translator:uav_burstcount
	signal nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata               : std_logic_vector(31 downto 0);  -- nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> nios2_qsys_grms_jtag_debug_module_translator:uav_writedata
	signal nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address                 : std_logic_vector(24 downto 0);  -- nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> nios2_qsys_grms_jtag_debug_module_translator:uav_address
	signal nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write                   : std_logic;                      -- nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> nios2_qsys_grms_jtag_debug_module_translator:uav_write
	signal nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock                    : std_logic;                      -- nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> nios2_qsys_grms_jtag_debug_module_translator:uav_lock
	signal nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read                    : std_logic;                      -- nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> nios2_qsys_grms_jtag_debug_module_translator:uav_read
	signal nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata                : std_logic_vector(31 downto 0);  -- nios2_qsys_grms_jtag_debug_module_translator:uav_readdata -> nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	signal nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid           : std_logic;                      -- nios2_qsys_grms_jtag_debug_module_translator:uav_readdatavalid -> nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess             : std_logic;                      -- nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> nios2_qsys_grms_jtag_debug_module_translator:uav_debugaccess
	signal nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable              : std_logic_vector(3 downto 0);   -- nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> nios2_qsys_grms_jtag_debug_module_translator:uav_byteenable
	signal nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket      : std_logic;                      -- nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid            : std_logic;                      -- nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket    : std_logic;                      -- nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data             : std_logic_vector(100 downto 0); -- nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready            : std_logic;                      -- nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket   : std_logic;                      -- nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid         : std_logic;                      -- nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket : std_logic;                      -- nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data          : std_logic_vector(100 downto 0); -- nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready         : std_logic;                      -- nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid       : std_logic;                      -- nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data        : std_logic_vector(33 downto 0);  -- nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready       : std_logic;                      -- nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest              : std_logic;                      -- jtag_uart_grms_avalon_jtag_slave_translator:uav_waitrequest -> jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount               : std_logic_vector(2 downto 0);   -- jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_uart_grms_avalon_jtag_slave_translator:uav_burstcount
	signal jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata                : std_logic_vector(31 downto 0);  -- jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_uart_grms_avalon_jtag_slave_translator:uav_writedata
	signal jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address                  : std_logic_vector(24 downto 0);  -- jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_uart_grms_avalon_jtag_slave_translator:uav_address
	signal jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write                    : std_logic;                      -- jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_uart_grms_avalon_jtag_slave_translator:uav_write
	signal jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock                     : std_logic;                      -- jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_uart_grms_avalon_jtag_slave_translator:uav_lock
	signal jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read                     : std_logic;                      -- jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_uart_grms_avalon_jtag_slave_translator:uav_read
	signal jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata                 : std_logic_vector(31 downto 0);  -- jtag_uart_grms_avalon_jtag_slave_translator:uav_readdata -> jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	signal jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid            : std_logic;                      -- jtag_uart_grms_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess              : std_logic;                      -- jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_uart_grms_avalon_jtag_slave_translator:uav_debugaccess
	signal jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable               : std_logic_vector(3 downto 0);   -- jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_uart_grms_avalon_jtag_slave_translator:uav_byteenable
	signal jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket       : std_logic;                      -- jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid             : std_logic;                      -- jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket     : std_logic;                      -- jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data              : std_logic_vector(100 downto 0); -- jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready             : std_logic;                      -- jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket    : std_logic;                      -- jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid          : std_logic;                      -- jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket  : std_logic;                      -- jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data           : std_logic_vector(100 downto 0); -- jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready          : std_logic;                      -- jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid        : std_logic;                      -- jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data         : std_logic_vector(33 downto 0);  -- jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready        : std_logic;                      -- jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                  : std_logic;                      -- new_sdram_controller_grms_s1_translator:uav_waitrequest -> new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                   : std_logic_vector(1 downto 0);   -- new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> new_sdram_controller_grms_s1_translator:uav_burstcount
	signal new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_m0_writedata                    : std_logic_vector(15 downto 0);  -- new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> new_sdram_controller_grms_s1_translator:uav_writedata
	signal new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_m0_address                      : std_logic_vector(24 downto 0);  -- new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent:m0_address -> new_sdram_controller_grms_s1_translator:uav_address
	signal new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_m0_write                        : std_logic;                      -- new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent:m0_write -> new_sdram_controller_grms_s1_translator:uav_write
	signal new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_m0_lock                         : std_logic;                      -- new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent:m0_lock -> new_sdram_controller_grms_s1_translator:uav_lock
	signal new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_m0_read                         : std_logic;                      -- new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent:m0_read -> new_sdram_controller_grms_s1_translator:uav_read
	signal new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_m0_readdata                     : std_logic_vector(15 downto 0);  -- new_sdram_controller_grms_s1_translator:uav_readdata -> new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                : std_logic;                      -- new_sdram_controller_grms_s1_translator:uav_readdatavalid -> new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                  : std_logic;                      -- new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> new_sdram_controller_grms_s1_translator:uav_debugaccess
	signal new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                   : std_logic_vector(1 downto 0);   -- new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> new_sdram_controller_grms_s1_translator:uav_byteenable
	signal new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket           : std_logic;                      -- new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                 : std_logic;                      -- new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket         : std_logic;                      -- new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_data                  : std_logic_vector(82 downto 0);  -- new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                 : std_logic;                      -- new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket        : std_logic;                      -- new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid              : std_logic;                      -- new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket      : std_logic;                      -- new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data               : std_logic_vector(82 downto 0);  -- new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready              : std_logic;                      -- new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid            : std_logic;                      -- new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	signal new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data             : std_logic_vector(17 downto 0);  -- new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	signal new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready            : std_logic;                      -- new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid            : std_logic;                      -- new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data             : std_logic_vector(17 downto 0);  -- new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready            : std_logic;                      -- new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	signal timer_grms_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                 : std_logic;                      -- timer_grms_s1_translator:uav_waitrequest -> timer_grms_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal timer_grms_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                  : std_logic_vector(2 downto 0);   -- timer_grms_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> timer_grms_s1_translator:uav_burstcount
	signal timer_grms_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                   : std_logic_vector(31 downto 0);  -- timer_grms_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> timer_grms_s1_translator:uav_writedata
	signal timer_grms_s1_translator_avalon_universal_slave_0_agent_m0_address                                     : std_logic_vector(24 downto 0);  -- timer_grms_s1_translator_avalon_universal_slave_0_agent:m0_address -> timer_grms_s1_translator:uav_address
	signal timer_grms_s1_translator_avalon_universal_slave_0_agent_m0_write                                       : std_logic;                      -- timer_grms_s1_translator_avalon_universal_slave_0_agent:m0_write -> timer_grms_s1_translator:uav_write
	signal timer_grms_s1_translator_avalon_universal_slave_0_agent_m0_lock                                        : std_logic;                      -- timer_grms_s1_translator_avalon_universal_slave_0_agent:m0_lock -> timer_grms_s1_translator:uav_lock
	signal timer_grms_s1_translator_avalon_universal_slave_0_agent_m0_read                                        : std_logic;                      -- timer_grms_s1_translator_avalon_universal_slave_0_agent:m0_read -> timer_grms_s1_translator:uav_read
	signal timer_grms_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                    : std_logic_vector(31 downto 0);  -- timer_grms_s1_translator:uav_readdata -> timer_grms_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal timer_grms_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                               : std_logic;                      -- timer_grms_s1_translator:uav_readdatavalid -> timer_grms_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal timer_grms_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                 : std_logic;                      -- timer_grms_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> timer_grms_s1_translator:uav_debugaccess
	signal timer_grms_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                  : std_logic_vector(3 downto 0);   -- timer_grms_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> timer_grms_s1_translator:uav_byteenable
	signal timer_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                          : std_logic;                      -- timer_grms_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> timer_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal timer_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                : std_logic;                      -- timer_grms_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> timer_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal timer_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                        : std_logic;                      -- timer_grms_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> timer_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal timer_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                 : std_logic_vector(100 downto 0); -- timer_grms_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> timer_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal timer_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                : std_logic;                      -- timer_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> timer_grms_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal timer_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                       : std_logic;                      -- timer_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> timer_grms_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal timer_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                             : std_logic;                      -- timer_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> timer_grms_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal timer_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                     : std_logic;                      -- timer_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> timer_grms_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal timer_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                              : std_logic_vector(100 downto 0); -- timer_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> timer_grms_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal timer_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                             : std_logic;                      -- timer_grms_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> timer_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal timer_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                           : std_logic;                      -- timer_grms_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> timer_grms_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal timer_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                            : std_logic_vector(33 downto 0);  -- timer_grms_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> timer_grms_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal timer_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                           : std_logic;                      -- timer_grms_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> timer_grms_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest                  : std_logic;                      -- lcd_16207_grms_control_slave_translator:uav_waitrequest -> lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount                   : std_logic_vector(2 downto 0);   -- lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> lcd_16207_grms_control_slave_translator:uav_burstcount
	signal lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata                    : std_logic_vector(31 downto 0);  -- lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> lcd_16207_grms_control_slave_translator:uav_writedata
	signal lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_m0_address                      : std_logic_vector(24 downto 0);  -- lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> lcd_16207_grms_control_slave_translator:uav_address
	signal lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_m0_write                        : std_logic;                      -- lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> lcd_16207_grms_control_slave_translator:uav_write
	signal lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_m0_lock                         : std_logic;                      -- lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> lcd_16207_grms_control_slave_translator:uav_lock
	signal lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_m0_read                         : std_logic;                      -- lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> lcd_16207_grms_control_slave_translator:uav_read
	signal lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata                     : std_logic_vector(31 downto 0);  -- lcd_16207_grms_control_slave_translator:uav_readdata -> lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	signal lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid                : std_logic;                      -- lcd_16207_grms_control_slave_translator:uav_readdatavalid -> lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess                  : std_logic;                      -- lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> lcd_16207_grms_control_slave_translator:uav_debugaccess
	signal lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable                   : std_logic_vector(3 downto 0);   -- lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> lcd_16207_grms_control_slave_translator:uav_byteenable
	signal lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket           : std_logic;                      -- lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid                 : std_logic;                      -- lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket         : std_logic;                      -- lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data                  : std_logic_vector(100 downto 0); -- lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready                 : std_logic;                      -- lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket        : std_logic;                      -- lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid              : std_logic;                      -- lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket      : std_logic;                      -- lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data               : std_logic_vector(100 downto 0); -- lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready              : std_logic;                      -- lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid            : std_logic;                      -- lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data             : std_logic_vector(33 downto 0);  -- lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready            : std_logic;                      -- lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal pa_grms_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                    : std_logic;                      -- pa_grms_s1_translator:uav_waitrequest -> pa_grms_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal pa_grms_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                     : std_logic_vector(2 downto 0);   -- pa_grms_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pa_grms_s1_translator:uav_burstcount
	signal pa_grms_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                      : std_logic_vector(31 downto 0);  -- pa_grms_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pa_grms_s1_translator:uav_writedata
	signal pa_grms_s1_translator_avalon_universal_slave_0_agent_m0_address                                        : std_logic_vector(24 downto 0);  -- pa_grms_s1_translator_avalon_universal_slave_0_agent:m0_address -> pa_grms_s1_translator:uav_address
	signal pa_grms_s1_translator_avalon_universal_slave_0_agent_m0_write                                          : std_logic;                      -- pa_grms_s1_translator_avalon_universal_slave_0_agent:m0_write -> pa_grms_s1_translator:uav_write
	signal pa_grms_s1_translator_avalon_universal_slave_0_agent_m0_lock                                           : std_logic;                      -- pa_grms_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pa_grms_s1_translator:uav_lock
	signal pa_grms_s1_translator_avalon_universal_slave_0_agent_m0_read                                           : std_logic;                      -- pa_grms_s1_translator_avalon_universal_slave_0_agent:m0_read -> pa_grms_s1_translator:uav_read
	signal pa_grms_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                       : std_logic_vector(31 downto 0);  -- pa_grms_s1_translator:uav_readdata -> pa_grms_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal pa_grms_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                  : std_logic;                      -- pa_grms_s1_translator:uav_readdatavalid -> pa_grms_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal pa_grms_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                    : std_logic;                      -- pa_grms_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pa_grms_s1_translator:uav_debugaccess
	signal pa_grms_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                     : std_logic_vector(3 downto 0);   -- pa_grms_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pa_grms_s1_translator:uav_byteenable
	signal pa_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                             : std_logic;                      -- pa_grms_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pa_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal pa_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                   : std_logic;                      -- pa_grms_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pa_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal pa_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                           : std_logic;                      -- pa_grms_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pa_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal pa_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                    : std_logic_vector(100 downto 0); -- pa_grms_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pa_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal pa_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                   : std_logic;                      -- pa_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pa_grms_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal pa_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                          : std_logic;                      -- pa_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pa_grms_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal pa_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                                : std_logic;                      -- pa_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pa_grms_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal pa_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                        : std_logic;                      -- pa_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pa_grms_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal pa_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                 : std_logic_vector(100 downto 0); -- pa_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pa_grms_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal pa_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                                : std_logic;                      -- pa_grms_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pa_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal pa_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                              : std_logic;                      -- pa_grms_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pa_grms_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal pa_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                               : std_logic_vector(33 downto 0);  -- pa_grms_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pa_grms_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal pa_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                              : std_logic;                      -- pa_grms_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pa_grms_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal pb_grms_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                    : std_logic;                      -- pb_grms_s1_translator:uav_waitrequest -> pb_grms_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal pb_grms_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                     : std_logic_vector(2 downto 0);   -- pb_grms_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pb_grms_s1_translator:uav_burstcount
	signal pb_grms_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                      : std_logic_vector(31 downto 0);  -- pb_grms_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pb_grms_s1_translator:uav_writedata
	signal pb_grms_s1_translator_avalon_universal_slave_0_agent_m0_address                                        : std_logic_vector(24 downto 0);  -- pb_grms_s1_translator_avalon_universal_slave_0_agent:m0_address -> pb_grms_s1_translator:uav_address
	signal pb_grms_s1_translator_avalon_universal_slave_0_agent_m0_write                                          : std_logic;                      -- pb_grms_s1_translator_avalon_universal_slave_0_agent:m0_write -> pb_grms_s1_translator:uav_write
	signal pb_grms_s1_translator_avalon_universal_slave_0_agent_m0_lock                                           : std_logic;                      -- pb_grms_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pb_grms_s1_translator:uav_lock
	signal pb_grms_s1_translator_avalon_universal_slave_0_agent_m0_read                                           : std_logic;                      -- pb_grms_s1_translator_avalon_universal_slave_0_agent:m0_read -> pb_grms_s1_translator:uav_read
	signal pb_grms_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                       : std_logic_vector(31 downto 0);  -- pb_grms_s1_translator:uav_readdata -> pb_grms_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal pb_grms_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                  : std_logic;                      -- pb_grms_s1_translator:uav_readdatavalid -> pb_grms_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal pb_grms_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                    : std_logic;                      -- pb_grms_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pb_grms_s1_translator:uav_debugaccess
	signal pb_grms_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                     : std_logic_vector(3 downto 0);   -- pb_grms_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pb_grms_s1_translator:uav_byteenable
	signal pb_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                             : std_logic;                      -- pb_grms_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pb_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal pb_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                   : std_logic;                      -- pb_grms_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pb_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal pb_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                           : std_logic;                      -- pb_grms_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pb_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal pb_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                    : std_logic_vector(100 downto 0); -- pb_grms_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pb_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal pb_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                   : std_logic;                      -- pb_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pb_grms_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal pb_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                          : std_logic;                      -- pb_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pb_grms_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal pb_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                                : std_logic;                      -- pb_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pb_grms_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal pb_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                        : std_logic;                      -- pb_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pb_grms_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal pb_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                 : std_logic_vector(100 downto 0); -- pb_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pb_grms_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal pb_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                                : std_logic;                      -- pb_grms_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pb_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal pb_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                              : std_logic;                      -- pb_grms_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pb_grms_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal pb_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                               : std_logic_vector(33 downto 0);  -- pb_grms_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pb_grms_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal pb_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                              : std_logic;                      -- pb_grms_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pb_grms_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal pc_grms_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                    : std_logic;                      -- pc_grms_s1_translator:uav_waitrequest -> pc_grms_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal pc_grms_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                     : std_logic_vector(2 downto 0);   -- pc_grms_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pc_grms_s1_translator:uav_burstcount
	signal pc_grms_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                      : std_logic_vector(31 downto 0);  -- pc_grms_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pc_grms_s1_translator:uav_writedata
	signal pc_grms_s1_translator_avalon_universal_slave_0_agent_m0_address                                        : std_logic_vector(24 downto 0);  -- pc_grms_s1_translator_avalon_universal_slave_0_agent:m0_address -> pc_grms_s1_translator:uav_address
	signal pc_grms_s1_translator_avalon_universal_slave_0_agent_m0_write                                          : std_logic;                      -- pc_grms_s1_translator_avalon_universal_slave_0_agent:m0_write -> pc_grms_s1_translator:uav_write
	signal pc_grms_s1_translator_avalon_universal_slave_0_agent_m0_lock                                           : std_logic;                      -- pc_grms_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pc_grms_s1_translator:uav_lock
	signal pc_grms_s1_translator_avalon_universal_slave_0_agent_m0_read                                           : std_logic;                      -- pc_grms_s1_translator_avalon_universal_slave_0_agent:m0_read -> pc_grms_s1_translator:uav_read
	signal pc_grms_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                       : std_logic_vector(31 downto 0);  -- pc_grms_s1_translator:uav_readdata -> pc_grms_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal pc_grms_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                  : std_logic;                      -- pc_grms_s1_translator:uav_readdatavalid -> pc_grms_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal pc_grms_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                    : std_logic;                      -- pc_grms_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pc_grms_s1_translator:uav_debugaccess
	signal pc_grms_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                     : std_logic_vector(3 downto 0);   -- pc_grms_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pc_grms_s1_translator:uav_byteenable
	signal pc_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                             : std_logic;                      -- pc_grms_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pc_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal pc_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                   : std_logic;                      -- pc_grms_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pc_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal pc_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                           : std_logic;                      -- pc_grms_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pc_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal pc_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                    : std_logic_vector(100 downto 0); -- pc_grms_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pc_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal pc_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                   : std_logic;                      -- pc_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pc_grms_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal pc_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                          : std_logic;                      -- pc_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pc_grms_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal pc_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                                : std_logic;                      -- pc_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pc_grms_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal pc_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                        : std_logic;                      -- pc_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pc_grms_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal pc_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                 : std_logic_vector(100 downto 0); -- pc_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pc_grms_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal pc_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                                : std_logic;                      -- pc_grms_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pc_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal pc_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                              : std_logic;                      -- pc_grms_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pc_grms_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal pc_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                               : std_logic_vector(33 downto 0);  -- pc_grms_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pc_grms_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal pc_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                              : std_logic;                      -- pc_grms_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pc_grms_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal pd_grms_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                    : std_logic;                      -- pd_grms_s1_translator:uav_waitrequest -> pd_grms_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal pd_grms_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                     : std_logic_vector(2 downto 0);   -- pd_grms_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pd_grms_s1_translator:uav_burstcount
	signal pd_grms_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                      : std_logic_vector(31 downto 0);  -- pd_grms_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pd_grms_s1_translator:uav_writedata
	signal pd_grms_s1_translator_avalon_universal_slave_0_agent_m0_address                                        : std_logic_vector(24 downto 0);  -- pd_grms_s1_translator_avalon_universal_slave_0_agent:m0_address -> pd_grms_s1_translator:uav_address
	signal pd_grms_s1_translator_avalon_universal_slave_0_agent_m0_write                                          : std_logic;                      -- pd_grms_s1_translator_avalon_universal_slave_0_agent:m0_write -> pd_grms_s1_translator:uav_write
	signal pd_grms_s1_translator_avalon_universal_slave_0_agent_m0_lock                                           : std_logic;                      -- pd_grms_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pd_grms_s1_translator:uav_lock
	signal pd_grms_s1_translator_avalon_universal_slave_0_agent_m0_read                                           : std_logic;                      -- pd_grms_s1_translator_avalon_universal_slave_0_agent:m0_read -> pd_grms_s1_translator:uav_read
	signal pd_grms_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                       : std_logic_vector(31 downto 0);  -- pd_grms_s1_translator:uav_readdata -> pd_grms_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal pd_grms_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                  : std_logic;                      -- pd_grms_s1_translator:uav_readdatavalid -> pd_grms_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal pd_grms_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                    : std_logic;                      -- pd_grms_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pd_grms_s1_translator:uav_debugaccess
	signal pd_grms_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                     : std_logic_vector(3 downto 0);   -- pd_grms_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pd_grms_s1_translator:uav_byteenable
	signal pd_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                             : std_logic;                      -- pd_grms_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pd_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal pd_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                   : std_logic;                      -- pd_grms_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pd_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal pd_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                           : std_logic;                      -- pd_grms_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pd_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal pd_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                    : std_logic_vector(100 downto 0); -- pd_grms_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pd_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal pd_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                   : std_logic;                      -- pd_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pd_grms_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal pd_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                          : std_logic;                      -- pd_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pd_grms_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal pd_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                                : std_logic;                      -- pd_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pd_grms_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal pd_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                        : std_logic;                      -- pd_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pd_grms_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal pd_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                 : std_logic_vector(100 downto 0); -- pd_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pd_grms_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal pd_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                                : std_logic;                      -- pd_grms_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pd_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal pd_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                              : std_logic;                      -- pd_grms_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pd_grms_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal pd_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                               : std_logic_vector(33 downto 0);  -- pd_grms_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pd_grms_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal pd_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                              : std_logic;                      -- pd_grms_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pd_grms_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal pe_grms_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                    : std_logic;                      -- pe_grms_s1_translator:uav_waitrequest -> pe_grms_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal pe_grms_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                     : std_logic_vector(2 downto 0);   -- pe_grms_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pe_grms_s1_translator:uav_burstcount
	signal pe_grms_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                      : std_logic_vector(31 downto 0);  -- pe_grms_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pe_grms_s1_translator:uav_writedata
	signal pe_grms_s1_translator_avalon_universal_slave_0_agent_m0_address                                        : std_logic_vector(24 downto 0);  -- pe_grms_s1_translator_avalon_universal_slave_0_agent:m0_address -> pe_grms_s1_translator:uav_address
	signal pe_grms_s1_translator_avalon_universal_slave_0_agent_m0_write                                          : std_logic;                      -- pe_grms_s1_translator_avalon_universal_slave_0_agent:m0_write -> pe_grms_s1_translator:uav_write
	signal pe_grms_s1_translator_avalon_universal_slave_0_agent_m0_lock                                           : std_logic;                      -- pe_grms_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pe_grms_s1_translator:uav_lock
	signal pe_grms_s1_translator_avalon_universal_slave_0_agent_m0_read                                           : std_logic;                      -- pe_grms_s1_translator_avalon_universal_slave_0_agent:m0_read -> pe_grms_s1_translator:uav_read
	signal pe_grms_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                       : std_logic_vector(31 downto 0);  -- pe_grms_s1_translator:uav_readdata -> pe_grms_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal pe_grms_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                  : std_logic;                      -- pe_grms_s1_translator:uav_readdatavalid -> pe_grms_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal pe_grms_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                    : std_logic;                      -- pe_grms_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pe_grms_s1_translator:uav_debugaccess
	signal pe_grms_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                     : std_logic_vector(3 downto 0);   -- pe_grms_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pe_grms_s1_translator:uav_byteenable
	signal pe_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                             : std_logic;                      -- pe_grms_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pe_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal pe_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                   : std_logic;                      -- pe_grms_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pe_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal pe_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                           : std_logic;                      -- pe_grms_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pe_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal pe_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                    : std_logic_vector(100 downto 0); -- pe_grms_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pe_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal pe_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                   : std_logic;                      -- pe_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pe_grms_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal pe_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                          : std_logic;                      -- pe_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pe_grms_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal pe_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                                : std_logic;                      -- pe_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pe_grms_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal pe_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                        : std_logic;                      -- pe_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pe_grms_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal pe_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                 : std_logic_vector(100 downto 0); -- pe_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pe_grms_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal pe_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                                : std_logic;                      -- pe_grms_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pe_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal pe_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                              : std_logic;                      -- pe_grms_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pe_grms_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal pe_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                               : std_logic_vector(33 downto 0);  -- pe_grms_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pe_grms_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal pe_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                              : std_logic;                      -- pe_grms_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pe_grms_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal pf_grms_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                    : std_logic;                      -- pf_grms_s1_translator:uav_waitrequest -> pf_grms_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal pf_grms_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                     : std_logic_vector(2 downto 0);   -- pf_grms_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pf_grms_s1_translator:uav_burstcount
	signal pf_grms_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                      : std_logic_vector(31 downto 0);  -- pf_grms_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pf_grms_s1_translator:uav_writedata
	signal pf_grms_s1_translator_avalon_universal_slave_0_agent_m0_address                                        : std_logic_vector(24 downto 0);  -- pf_grms_s1_translator_avalon_universal_slave_0_agent:m0_address -> pf_grms_s1_translator:uav_address
	signal pf_grms_s1_translator_avalon_universal_slave_0_agent_m0_write                                          : std_logic;                      -- pf_grms_s1_translator_avalon_universal_slave_0_agent:m0_write -> pf_grms_s1_translator:uav_write
	signal pf_grms_s1_translator_avalon_universal_slave_0_agent_m0_lock                                           : std_logic;                      -- pf_grms_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pf_grms_s1_translator:uav_lock
	signal pf_grms_s1_translator_avalon_universal_slave_0_agent_m0_read                                           : std_logic;                      -- pf_grms_s1_translator_avalon_universal_slave_0_agent:m0_read -> pf_grms_s1_translator:uav_read
	signal pf_grms_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                       : std_logic_vector(31 downto 0);  -- pf_grms_s1_translator:uav_readdata -> pf_grms_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal pf_grms_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                  : std_logic;                      -- pf_grms_s1_translator:uav_readdatavalid -> pf_grms_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal pf_grms_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                    : std_logic;                      -- pf_grms_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pf_grms_s1_translator:uav_debugaccess
	signal pf_grms_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                     : std_logic_vector(3 downto 0);   -- pf_grms_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pf_grms_s1_translator:uav_byteenable
	signal pf_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                             : std_logic;                      -- pf_grms_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pf_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal pf_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                   : std_logic;                      -- pf_grms_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pf_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal pf_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                           : std_logic;                      -- pf_grms_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pf_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal pf_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                    : std_logic_vector(100 downto 0); -- pf_grms_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pf_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal pf_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                   : std_logic;                      -- pf_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pf_grms_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal pf_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                          : std_logic;                      -- pf_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pf_grms_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal pf_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                                : std_logic;                      -- pf_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pf_grms_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal pf_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                        : std_logic;                      -- pf_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pf_grms_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal pf_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                 : std_logic_vector(100 downto 0); -- pf_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pf_grms_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal pf_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                                : std_logic;                      -- pf_grms_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pf_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal pf_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                              : std_logic;                      -- pf_grms_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pf_grms_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal pf_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                               : std_logic_vector(33 downto 0);  -- pf_grms_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pf_grms_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal pf_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                              : std_logic;                      -- pf_grms_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pf_grms_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal pg_grms_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                    : std_logic;                      -- pg_grms_s1_translator:uav_waitrequest -> pg_grms_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal pg_grms_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                     : std_logic_vector(2 downto 0);   -- pg_grms_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pg_grms_s1_translator:uav_burstcount
	signal pg_grms_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                      : std_logic_vector(31 downto 0);  -- pg_grms_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pg_grms_s1_translator:uav_writedata
	signal pg_grms_s1_translator_avalon_universal_slave_0_agent_m0_address                                        : std_logic_vector(24 downto 0);  -- pg_grms_s1_translator_avalon_universal_slave_0_agent:m0_address -> pg_grms_s1_translator:uav_address
	signal pg_grms_s1_translator_avalon_universal_slave_0_agent_m0_write                                          : std_logic;                      -- pg_grms_s1_translator_avalon_universal_slave_0_agent:m0_write -> pg_grms_s1_translator:uav_write
	signal pg_grms_s1_translator_avalon_universal_slave_0_agent_m0_lock                                           : std_logic;                      -- pg_grms_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pg_grms_s1_translator:uav_lock
	signal pg_grms_s1_translator_avalon_universal_slave_0_agent_m0_read                                           : std_logic;                      -- pg_grms_s1_translator_avalon_universal_slave_0_agent:m0_read -> pg_grms_s1_translator:uav_read
	signal pg_grms_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                       : std_logic_vector(31 downto 0);  -- pg_grms_s1_translator:uav_readdata -> pg_grms_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal pg_grms_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                  : std_logic;                      -- pg_grms_s1_translator:uav_readdatavalid -> pg_grms_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal pg_grms_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                    : std_logic;                      -- pg_grms_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pg_grms_s1_translator:uav_debugaccess
	signal pg_grms_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                     : std_logic_vector(3 downto 0);   -- pg_grms_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pg_grms_s1_translator:uav_byteenable
	signal pg_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                             : std_logic;                      -- pg_grms_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pg_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal pg_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                   : std_logic;                      -- pg_grms_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pg_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal pg_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                           : std_logic;                      -- pg_grms_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pg_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal pg_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                    : std_logic_vector(100 downto 0); -- pg_grms_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pg_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal pg_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                   : std_logic;                      -- pg_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pg_grms_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal pg_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                          : std_logic;                      -- pg_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pg_grms_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal pg_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                                : std_logic;                      -- pg_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pg_grms_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal pg_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                        : std_logic;                      -- pg_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pg_grms_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal pg_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                 : std_logic_vector(100 downto 0); -- pg_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pg_grms_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal pg_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                                : std_logic;                      -- pg_grms_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pg_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal pg_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                              : std_logic;                      -- pg_grms_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pg_grms_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal pg_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                               : std_logic_vector(33 downto 0);  -- pg_grms_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pg_grms_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal pg_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                              : std_logic;                      -- pg_grms_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pg_grms_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal ph_grms_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                    : std_logic;                      -- ph_grms_s1_translator:uav_waitrequest -> ph_grms_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal ph_grms_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                     : std_logic_vector(2 downto 0);   -- ph_grms_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> ph_grms_s1_translator:uav_burstcount
	signal ph_grms_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                      : std_logic_vector(31 downto 0);  -- ph_grms_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> ph_grms_s1_translator:uav_writedata
	signal ph_grms_s1_translator_avalon_universal_slave_0_agent_m0_address                                        : std_logic_vector(24 downto 0);  -- ph_grms_s1_translator_avalon_universal_slave_0_agent:m0_address -> ph_grms_s1_translator:uav_address
	signal ph_grms_s1_translator_avalon_universal_slave_0_agent_m0_write                                          : std_logic;                      -- ph_grms_s1_translator_avalon_universal_slave_0_agent:m0_write -> ph_grms_s1_translator:uav_write
	signal ph_grms_s1_translator_avalon_universal_slave_0_agent_m0_lock                                           : std_logic;                      -- ph_grms_s1_translator_avalon_universal_slave_0_agent:m0_lock -> ph_grms_s1_translator:uav_lock
	signal ph_grms_s1_translator_avalon_universal_slave_0_agent_m0_read                                           : std_logic;                      -- ph_grms_s1_translator_avalon_universal_slave_0_agent:m0_read -> ph_grms_s1_translator:uav_read
	signal ph_grms_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                       : std_logic_vector(31 downto 0);  -- ph_grms_s1_translator:uav_readdata -> ph_grms_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal ph_grms_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                  : std_logic;                      -- ph_grms_s1_translator:uav_readdatavalid -> ph_grms_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal ph_grms_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                    : std_logic;                      -- ph_grms_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> ph_grms_s1_translator:uav_debugaccess
	signal ph_grms_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                     : std_logic_vector(3 downto 0);   -- ph_grms_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> ph_grms_s1_translator:uav_byteenable
	signal ph_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                             : std_logic;                      -- ph_grms_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> ph_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal ph_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                   : std_logic;                      -- ph_grms_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> ph_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal ph_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                           : std_logic;                      -- ph_grms_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> ph_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal ph_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                    : std_logic_vector(100 downto 0); -- ph_grms_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> ph_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal ph_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                   : std_logic;                      -- ph_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> ph_grms_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal ph_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                          : std_logic;                      -- ph_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> ph_grms_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal ph_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                                : std_logic;                      -- ph_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> ph_grms_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal ph_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                        : std_logic;                      -- ph_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> ph_grms_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal ph_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                 : std_logic_vector(100 downto 0); -- ph_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> ph_grms_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal ph_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                                : std_logic;                      -- ph_grms_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> ph_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal ph_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                              : std_logic;                      -- ph_grms_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> ph_grms_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal ph_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                               : std_logic_vector(33 downto 0);  -- ph_grms_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> ph_grms_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal ph_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                              : std_logic;                      -- ph_grms_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> ph_grms_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal pi_grms_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                    : std_logic;                      -- pi_grms_s1_translator:uav_waitrequest -> pi_grms_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal pi_grms_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                     : std_logic_vector(2 downto 0);   -- pi_grms_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pi_grms_s1_translator:uav_burstcount
	signal pi_grms_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                      : std_logic_vector(31 downto 0);  -- pi_grms_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pi_grms_s1_translator:uav_writedata
	signal pi_grms_s1_translator_avalon_universal_slave_0_agent_m0_address                                        : std_logic_vector(24 downto 0);  -- pi_grms_s1_translator_avalon_universal_slave_0_agent:m0_address -> pi_grms_s1_translator:uav_address
	signal pi_grms_s1_translator_avalon_universal_slave_0_agent_m0_write                                          : std_logic;                      -- pi_grms_s1_translator_avalon_universal_slave_0_agent:m0_write -> pi_grms_s1_translator:uav_write
	signal pi_grms_s1_translator_avalon_universal_slave_0_agent_m0_lock                                           : std_logic;                      -- pi_grms_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pi_grms_s1_translator:uav_lock
	signal pi_grms_s1_translator_avalon_universal_slave_0_agent_m0_read                                           : std_logic;                      -- pi_grms_s1_translator_avalon_universal_slave_0_agent:m0_read -> pi_grms_s1_translator:uav_read
	signal pi_grms_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                       : std_logic_vector(31 downto 0);  -- pi_grms_s1_translator:uav_readdata -> pi_grms_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal pi_grms_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                  : std_logic;                      -- pi_grms_s1_translator:uav_readdatavalid -> pi_grms_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal pi_grms_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                    : std_logic;                      -- pi_grms_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pi_grms_s1_translator:uav_debugaccess
	signal pi_grms_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                     : std_logic_vector(3 downto 0);   -- pi_grms_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pi_grms_s1_translator:uav_byteenable
	signal pi_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                             : std_logic;                      -- pi_grms_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pi_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal pi_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                   : std_logic;                      -- pi_grms_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pi_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal pi_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                           : std_logic;                      -- pi_grms_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pi_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal pi_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                    : std_logic_vector(100 downto 0); -- pi_grms_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pi_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal pi_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                   : std_logic;                      -- pi_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pi_grms_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal pi_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                          : std_logic;                      -- pi_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pi_grms_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal pi_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                                : std_logic;                      -- pi_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pi_grms_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal pi_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                        : std_logic;                      -- pi_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pi_grms_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal pi_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                 : std_logic_vector(100 downto 0); -- pi_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pi_grms_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal pi_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                                : std_logic;                      -- pi_grms_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pi_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal pi_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                              : std_logic;                      -- pi_grms_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pi_grms_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal pi_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                               : std_logic_vector(33 downto 0);  -- pi_grms_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pi_grms_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal pi_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                              : std_logic;                      -- pi_grms_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pi_grms_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal nios2_qsys_grms_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket           : std_logic;                      -- nios2_qsys_grms_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	signal nios2_qsys_grms_instruction_master_translator_avalon_universal_master_0_agent_cp_valid                 : std_logic;                      -- nios2_qsys_grms_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	signal nios2_qsys_grms_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket         : std_logic;                      -- nios2_qsys_grms_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	signal nios2_qsys_grms_instruction_master_translator_avalon_universal_master_0_agent_cp_data                  : std_logic_vector(99 downto 0);  -- nios2_qsys_grms_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	signal nios2_qsys_grms_instruction_master_translator_avalon_universal_master_0_agent_cp_ready                 : std_logic;                      -- addr_router:sink_ready -> nios2_qsys_grms_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	signal nios2_qsys_grms_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket                  : std_logic;                      -- nios2_qsys_grms_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	signal nios2_qsys_grms_data_master_translator_avalon_universal_master_0_agent_cp_valid                        : std_logic;                      -- nios2_qsys_grms_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	signal nios2_qsys_grms_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket                : std_logic;                      -- nios2_qsys_grms_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	signal nios2_qsys_grms_data_master_translator_avalon_universal_master_0_agent_cp_data                         : std_logic_vector(99 downto 0);  -- nios2_qsys_grms_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	signal nios2_qsys_grms_data_master_translator_avalon_universal_master_0_agent_cp_ready                        : std_logic;                      -- addr_router_001:sink_ready -> nios2_qsys_grms_data_master_translator_avalon_universal_master_0_agent:cp_ready
	signal nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket             : std_logic;                      -- nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	signal nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid                   : std_logic;                      -- nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	signal nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket           : std_logic;                      -- nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	signal nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data                    : std_logic_vector(99 downto 0);  -- nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	signal nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready                   : std_logic;                      -- id_router:sink_ready -> nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	signal jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket              : std_logic;                      -- jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	signal jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid                    : std_logic;                      -- jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	signal jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket            : std_logic;                      -- jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	signal jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data                     : std_logic_vector(99 downto 0);  -- jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	signal jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready                    : std_logic;                      -- id_router_001:sink_ready -> jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	signal new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                  : std_logic;                      -- new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	signal new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rp_valid                        : std_logic;                      -- new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	signal new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                : std_logic;                      -- new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	signal new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rp_data                         : std_logic_vector(81 downto 0);  -- new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	signal new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rp_ready                        : std_logic;                      -- id_router_002:sink_ready -> new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal timer_grms_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                 : std_logic;                      -- timer_grms_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	signal timer_grms_s1_translator_avalon_universal_slave_0_agent_rp_valid                                       : std_logic;                      -- timer_grms_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	signal timer_grms_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                               : std_logic;                      -- timer_grms_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	signal timer_grms_s1_translator_avalon_universal_slave_0_agent_rp_data                                        : std_logic_vector(99 downto 0);  -- timer_grms_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	signal timer_grms_s1_translator_avalon_universal_slave_0_agent_rp_ready                                       : std_logic;                      -- id_router_003:sink_ready -> timer_grms_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket                  : std_logic;                      -- lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	signal lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_rp_valid                        : std_logic;                      -- lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	signal lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket                : std_logic;                      -- lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	signal lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_rp_data                         : std_logic_vector(99 downto 0);  -- lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	signal lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_rp_ready                        : std_logic;                      -- id_router_004:sink_ready -> lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	signal pa_grms_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                    : std_logic;                      -- pa_grms_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	signal pa_grms_s1_translator_avalon_universal_slave_0_agent_rp_valid                                          : std_logic;                      -- pa_grms_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	signal pa_grms_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                  : std_logic;                      -- pa_grms_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	signal pa_grms_s1_translator_avalon_universal_slave_0_agent_rp_data                                           : std_logic_vector(99 downto 0);  -- pa_grms_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	signal pa_grms_s1_translator_avalon_universal_slave_0_agent_rp_ready                                          : std_logic;                      -- id_router_005:sink_ready -> pa_grms_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal pb_grms_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                    : std_logic;                      -- pb_grms_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	signal pb_grms_s1_translator_avalon_universal_slave_0_agent_rp_valid                                          : std_logic;                      -- pb_grms_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	signal pb_grms_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                  : std_logic;                      -- pb_grms_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	signal pb_grms_s1_translator_avalon_universal_slave_0_agent_rp_data                                           : std_logic_vector(99 downto 0);  -- pb_grms_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	signal pb_grms_s1_translator_avalon_universal_slave_0_agent_rp_ready                                          : std_logic;                      -- id_router_006:sink_ready -> pb_grms_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal pc_grms_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                    : std_logic;                      -- pc_grms_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_007:sink_endofpacket
	signal pc_grms_s1_translator_avalon_universal_slave_0_agent_rp_valid                                          : std_logic;                      -- pc_grms_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_007:sink_valid
	signal pc_grms_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                  : std_logic;                      -- pc_grms_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_007:sink_startofpacket
	signal pc_grms_s1_translator_avalon_universal_slave_0_agent_rp_data                                           : std_logic_vector(99 downto 0);  -- pc_grms_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_007:sink_data
	signal pc_grms_s1_translator_avalon_universal_slave_0_agent_rp_ready                                          : std_logic;                      -- id_router_007:sink_ready -> pc_grms_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal pd_grms_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                    : std_logic;                      -- pd_grms_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_008:sink_endofpacket
	signal pd_grms_s1_translator_avalon_universal_slave_0_agent_rp_valid                                          : std_logic;                      -- pd_grms_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_008:sink_valid
	signal pd_grms_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                  : std_logic;                      -- pd_grms_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_008:sink_startofpacket
	signal pd_grms_s1_translator_avalon_universal_slave_0_agent_rp_data                                           : std_logic_vector(99 downto 0);  -- pd_grms_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_008:sink_data
	signal pd_grms_s1_translator_avalon_universal_slave_0_agent_rp_ready                                          : std_logic;                      -- id_router_008:sink_ready -> pd_grms_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal pe_grms_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                    : std_logic;                      -- pe_grms_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_009:sink_endofpacket
	signal pe_grms_s1_translator_avalon_universal_slave_0_agent_rp_valid                                          : std_logic;                      -- pe_grms_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_009:sink_valid
	signal pe_grms_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                  : std_logic;                      -- pe_grms_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_009:sink_startofpacket
	signal pe_grms_s1_translator_avalon_universal_slave_0_agent_rp_data                                           : std_logic_vector(99 downto 0);  -- pe_grms_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_009:sink_data
	signal pe_grms_s1_translator_avalon_universal_slave_0_agent_rp_ready                                          : std_logic;                      -- id_router_009:sink_ready -> pe_grms_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal pf_grms_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                    : std_logic;                      -- pf_grms_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_010:sink_endofpacket
	signal pf_grms_s1_translator_avalon_universal_slave_0_agent_rp_valid                                          : std_logic;                      -- pf_grms_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_010:sink_valid
	signal pf_grms_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                  : std_logic;                      -- pf_grms_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_010:sink_startofpacket
	signal pf_grms_s1_translator_avalon_universal_slave_0_agent_rp_data                                           : std_logic_vector(99 downto 0);  -- pf_grms_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_010:sink_data
	signal pf_grms_s1_translator_avalon_universal_slave_0_agent_rp_ready                                          : std_logic;                      -- id_router_010:sink_ready -> pf_grms_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal pg_grms_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                    : std_logic;                      -- pg_grms_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_011:sink_endofpacket
	signal pg_grms_s1_translator_avalon_universal_slave_0_agent_rp_valid                                          : std_logic;                      -- pg_grms_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_011:sink_valid
	signal pg_grms_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                  : std_logic;                      -- pg_grms_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_011:sink_startofpacket
	signal pg_grms_s1_translator_avalon_universal_slave_0_agent_rp_data                                           : std_logic_vector(99 downto 0);  -- pg_grms_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_011:sink_data
	signal pg_grms_s1_translator_avalon_universal_slave_0_agent_rp_ready                                          : std_logic;                      -- id_router_011:sink_ready -> pg_grms_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal ph_grms_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                    : std_logic;                      -- ph_grms_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_012:sink_endofpacket
	signal ph_grms_s1_translator_avalon_universal_slave_0_agent_rp_valid                                          : std_logic;                      -- ph_grms_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_012:sink_valid
	signal ph_grms_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                  : std_logic;                      -- ph_grms_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_012:sink_startofpacket
	signal ph_grms_s1_translator_avalon_universal_slave_0_agent_rp_data                                           : std_logic_vector(99 downto 0);  -- ph_grms_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_012:sink_data
	signal ph_grms_s1_translator_avalon_universal_slave_0_agent_rp_ready                                          : std_logic;                      -- id_router_012:sink_ready -> ph_grms_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal pi_grms_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                    : std_logic;                      -- pi_grms_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_013:sink_endofpacket
	signal pi_grms_s1_translator_avalon_universal_slave_0_agent_rp_valid                                          : std_logic;                      -- pi_grms_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_013:sink_valid
	signal pi_grms_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                  : std_logic;                      -- pi_grms_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_013:sink_startofpacket
	signal pi_grms_s1_translator_avalon_universal_slave_0_agent_rp_data                                           : std_logic_vector(99 downto 0);  -- pi_grms_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_013:sink_data
	signal pi_grms_s1_translator_avalon_universal_slave_0_agent_rp_ready                                          : std_logic;                      -- id_router_013:sink_ready -> pi_grms_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal burst_adapter_source0_endofpacket                                                                      : std_logic;                      -- burst_adapter:source0_endofpacket -> new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal burst_adapter_source0_valid                                                                            : std_logic;                      -- burst_adapter:source0_valid -> new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal burst_adapter_source0_startofpacket                                                                    : std_logic;                      -- burst_adapter:source0_startofpacket -> new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal burst_adapter_source0_data                                                                             : std_logic_vector(81 downto 0);  -- burst_adapter:source0_data -> new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal burst_adapter_source0_ready                                                                            : std_logic;                      -- new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter:source0_ready
	signal burst_adapter_source0_channel                                                                          : std_logic_vector(13 downto 0);  -- burst_adapter:source0_channel -> new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal rst_controller_reset_out_reset                                                                         : std_logic;                      -- rst_controller:reset_out -> [addr_router:reset, addr_router_001:reset, burst_adapter:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_mux:reset, cmd_xbar_mux_001:reset, cmd_xbar_mux_002:reset, cmd_xbar_mux_003:reset, cmd_xbar_mux_004:reset, cmd_xbar_mux_005:reset, cmd_xbar_mux_006:reset, cmd_xbar_mux_007:reset, cmd_xbar_mux_008:reset, cmd_xbar_mux_009:reset, cmd_xbar_mux_010:reset, cmd_xbar_mux_011:reset, cmd_xbar_mux_012:reset, cmd_xbar_mux_013:reset, id_router:reset, id_router_001:reset, id_router_002:reset, id_router_003:reset, id_router_004:reset, id_router_005:reset, id_router_006:reset, id_router_007:reset, id_router_008:reset, id_router_009:reset, id_router_010:reset, id_router_011:reset, id_router_012:reset, id_router_013:reset, irq_mapper:reset, jtag_uart_grms_avalon_jtag_slave_translator:reset, jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, lcd_16207_grms_control_slave_translator:reset, lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent:reset, lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, new_sdram_controller_grms_s1_translator:reset, new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent:reset, new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, nios2_qsys_grms_data_master_translator:reset, nios2_qsys_grms_data_master_translator_avalon_universal_master_0_agent:reset, nios2_qsys_grms_instruction_master_translator:reset, nios2_qsys_grms_instruction_master_translator_avalon_universal_master_0_agent:reset, nios2_qsys_grms_jtag_debug_module_translator:reset, nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pa_grms_s1_translator:reset, pa_grms_s1_translator_avalon_universal_slave_0_agent:reset, pa_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pb_grms_s1_translator:reset, pb_grms_s1_translator_avalon_universal_slave_0_agent:reset, pb_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pc_grms_s1_translator:reset, pc_grms_s1_translator_avalon_universal_slave_0_agent:reset, pc_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pd_grms_s1_translator:reset, pd_grms_s1_translator_avalon_universal_slave_0_agent:reset, pd_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pe_grms_s1_translator:reset, pe_grms_s1_translator_avalon_universal_slave_0_agent:reset, pe_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pf_grms_s1_translator:reset, pf_grms_s1_translator_avalon_universal_slave_0_agent:reset, pf_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pg_grms_s1_translator:reset, pg_grms_s1_translator_avalon_universal_slave_0_agent:reset, pg_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, ph_grms_s1_translator:reset, ph_grms_s1_translator_avalon_universal_slave_0_agent:reset, ph_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pi_grms_s1_translator:reset, pi_grms_s1_translator_avalon_universal_slave_0_agent:reset, pi_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_004:reset, rsp_xbar_demux_005:reset, rsp_xbar_demux_006:reset, rsp_xbar_demux_007:reset, rsp_xbar_demux_008:reset, rsp_xbar_demux_009:reset, rsp_xbar_demux_010:reset, rsp_xbar_demux_011:reset, rsp_xbar_demux_012:reset, rsp_xbar_demux_013:reset, rsp_xbar_mux:reset, rsp_xbar_mux_001:reset, rst_controller_reset_out_reset:in, timer_grms_s1_translator:reset, timer_grms_s1_translator_avalon_universal_slave_0_agent:reset, timer_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, width_adapter:reset, width_adapter_001:reset]
	signal cmd_xbar_demux_src0_endofpacket                                                                        : std_logic;                      -- cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	signal cmd_xbar_demux_src0_valid                                                                              : std_logic;                      -- cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	signal cmd_xbar_demux_src0_startofpacket                                                                      : std_logic;                      -- cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	signal cmd_xbar_demux_src0_data                                                                               : std_logic_vector(99 downto 0);  -- cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	signal cmd_xbar_demux_src0_channel                                                                            : std_logic_vector(13 downto 0);  -- cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	signal cmd_xbar_demux_src0_ready                                                                              : std_logic;                      -- cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	signal cmd_xbar_demux_src1_endofpacket                                                                        : std_logic;                      -- cmd_xbar_demux:src1_endofpacket -> cmd_xbar_mux_001:sink0_endofpacket
	signal cmd_xbar_demux_src1_valid                                                                              : std_logic;                      -- cmd_xbar_demux:src1_valid -> cmd_xbar_mux_001:sink0_valid
	signal cmd_xbar_demux_src1_startofpacket                                                                      : std_logic;                      -- cmd_xbar_demux:src1_startofpacket -> cmd_xbar_mux_001:sink0_startofpacket
	signal cmd_xbar_demux_src1_data                                                                               : std_logic_vector(99 downto 0);  -- cmd_xbar_demux:src1_data -> cmd_xbar_mux_001:sink0_data
	signal cmd_xbar_demux_src1_channel                                                                            : std_logic_vector(13 downto 0);  -- cmd_xbar_demux:src1_channel -> cmd_xbar_mux_001:sink0_channel
	signal cmd_xbar_demux_src1_ready                                                                              : std_logic;                      -- cmd_xbar_mux_001:sink0_ready -> cmd_xbar_demux:src1_ready
	signal cmd_xbar_demux_src2_endofpacket                                                                        : std_logic;                      -- cmd_xbar_demux:src2_endofpacket -> cmd_xbar_mux_002:sink0_endofpacket
	signal cmd_xbar_demux_src2_valid                                                                              : std_logic;                      -- cmd_xbar_demux:src2_valid -> cmd_xbar_mux_002:sink0_valid
	signal cmd_xbar_demux_src2_startofpacket                                                                      : std_logic;                      -- cmd_xbar_demux:src2_startofpacket -> cmd_xbar_mux_002:sink0_startofpacket
	signal cmd_xbar_demux_src2_data                                                                               : std_logic_vector(99 downto 0);  -- cmd_xbar_demux:src2_data -> cmd_xbar_mux_002:sink0_data
	signal cmd_xbar_demux_src2_channel                                                                            : std_logic_vector(13 downto 0);  -- cmd_xbar_demux:src2_channel -> cmd_xbar_mux_002:sink0_channel
	signal cmd_xbar_demux_src2_ready                                                                              : std_logic;                      -- cmd_xbar_mux_002:sink0_ready -> cmd_xbar_demux:src2_ready
	signal cmd_xbar_demux_src3_endofpacket                                                                        : std_logic;                      -- cmd_xbar_demux:src3_endofpacket -> cmd_xbar_mux_003:sink0_endofpacket
	signal cmd_xbar_demux_src3_valid                                                                              : std_logic;                      -- cmd_xbar_demux:src3_valid -> cmd_xbar_mux_003:sink0_valid
	signal cmd_xbar_demux_src3_startofpacket                                                                      : std_logic;                      -- cmd_xbar_demux:src3_startofpacket -> cmd_xbar_mux_003:sink0_startofpacket
	signal cmd_xbar_demux_src3_data                                                                               : std_logic_vector(99 downto 0);  -- cmd_xbar_demux:src3_data -> cmd_xbar_mux_003:sink0_data
	signal cmd_xbar_demux_src3_channel                                                                            : std_logic_vector(13 downto 0);  -- cmd_xbar_demux:src3_channel -> cmd_xbar_mux_003:sink0_channel
	signal cmd_xbar_demux_src3_ready                                                                              : std_logic;                      -- cmd_xbar_mux_003:sink0_ready -> cmd_xbar_demux:src3_ready
	signal cmd_xbar_demux_src4_endofpacket                                                                        : std_logic;                      -- cmd_xbar_demux:src4_endofpacket -> cmd_xbar_mux_004:sink0_endofpacket
	signal cmd_xbar_demux_src4_valid                                                                              : std_logic;                      -- cmd_xbar_demux:src4_valid -> cmd_xbar_mux_004:sink0_valid
	signal cmd_xbar_demux_src4_startofpacket                                                                      : std_logic;                      -- cmd_xbar_demux:src4_startofpacket -> cmd_xbar_mux_004:sink0_startofpacket
	signal cmd_xbar_demux_src4_data                                                                               : std_logic_vector(99 downto 0);  -- cmd_xbar_demux:src4_data -> cmd_xbar_mux_004:sink0_data
	signal cmd_xbar_demux_src4_channel                                                                            : std_logic_vector(13 downto 0);  -- cmd_xbar_demux:src4_channel -> cmd_xbar_mux_004:sink0_channel
	signal cmd_xbar_demux_src4_ready                                                                              : std_logic;                      -- cmd_xbar_mux_004:sink0_ready -> cmd_xbar_demux:src4_ready
	signal cmd_xbar_demux_src5_endofpacket                                                                        : std_logic;                      -- cmd_xbar_demux:src5_endofpacket -> cmd_xbar_mux_005:sink0_endofpacket
	signal cmd_xbar_demux_src5_valid                                                                              : std_logic;                      -- cmd_xbar_demux:src5_valid -> cmd_xbar_mux_005:sink0_valid
	signal cmd_xbar_demux_src5_startofpacket                                                                      : std_logic;                      -- cmd_xbar_demux:src5_startofpacket -> cmd_xbar_mux_005:sink0_startofpacket
	signal cmd_xbar_demux_src5_data                                                                               : std_logic_vector(99 downto 0);  -- cmd_xbar_demux:src5_data -> cmd_xbar_mux_005:sink0_data
	signal cmd_xbar_demux_src5_channel                                                                            : std_logic_vector(13 downto 0);  -- cmd_xbar_demux:src5_channel -> cmd_xbar_mux_005:sink0_channel
	signal cmd_xbar_demux_src5_ready                                                                              : std_logic;                      -- cmd_xbar_mux_005:sink0_ready -> cmd_xbar_demux:src5_ready
	signal cmd_xbar_demux_src6_endofpacket                                                                        : std_logic;                      -- cmd_xbar_demux:src6_endofpacket -> cmd_xbar_mux_006:sink0_endofpacket
	signal cmd_xbar_demux_src6_valid                                                                              : std_logic;                      -- cmd_xbar_demux:src6_valid -> cmd_xbar_mux_006:sink0_valid
	signal cmd_xbar_demux_src6_startofpacket                                                                      : std_logic;                      -- cmd_xbar_demux:src6_startofpacket -> cmd_xbar_mux_006:sink0_startofpacket
	signal cmd_xbar_demux_src6_data                                                                               : std_logic_vector(99 downto 0);  -- cmd_xbar_demux:src6_data -> cmd_xbar_mux_006:sink0_data
	signal cmd_xbar_demux_src6_channel                                                                            : std_logic_vector(13 downto 0);  -- cmd_xbar_demux:src6_channel -> cmd_xbar_mux_006:sink0_channel
	signal cmd_xbar_demux_src6_ready                                                                              : std_logic;                      -- cmd_xbar_mux_006:sink0_ready -> cmd_xbar_demux:src6_ready
	signal cmd_xbar_demux_src7_endofpacket                                                                        : std_logic;                      -- cmd_xbar_demux:src7_endofpacket -> cmd_xbar_mux_007:sink0_endofpacket
	signal cmd_xbar_demux_src7_valid                                                                              : std_logic;                      -- cmd_xbar_demux:src7_valid -> cmd_xbar_mux_007:sink0_valid
	signal cmd_xbar_demux_src7_startofpacket                                                                      : std_logic;                      -- cmd_xbar_demux:src7_startofpacket -> cmd_xbar_mux_007:sink0_startofpacket
	signal cmd_xbar_demux_src7_data                                                                               : std_logic_vector(99 downto 0);  -- cmd_xbar_demux:src7_data -> cmd_xbar_mux_007:sink0_data
	signal cmd_xbar_demux_src7_channel                                                                            : std_logic_vector(13 downto 0);  -- cmd_xbar_demux:src7_channel -> cmd_xbar_mux_007:sink0_channel
	signal cmd_xbar_demux_src7_ready                                                                              : std_logic;                      -- cmd_xbar_mux_007:sink0_ready -> cmd_xbar_demux:src7_ready
	signal cmd_xbar_demux_src8_endofpacket                                                                        : std_logic;                      -- cmd_xbar_demux:src8_endofpacket -> cmd_xbar_mux_008:sink0_endofpacket
	signal cmd_xbar_demux_src8_valid                                                                              : std_logic;                      -- cmd_xbar_demux:src8_valid -> cmd_xbar_mux_008:sink0_valid
	signal cmd_xbar_demux_src8_startofpacket                                                                      : std_logic;                      -- cmd_xbar_demux:src8_startofpacket -> cmd_xbar_mux_008:sink0_startofpacket
	signal cmd_xbar_demux_src8_data                                                                               : std_logic_vector(99 downto 0);  -- cmd_xbar_demux:src8_data -> cmd_xbar_mux_008:sink0_data
	signal cmd_xbar_demux_src8_channel                                                                            : std_logic_vector(13 downto 0);  -- cmd_xbar_demux:src8_channel -> cmd_xbar_mux_008:sink0_channel
	signal cmd_xbar_demux_src8_ready                                                                              : std_logic;                      -- cmd_xbar_mux_008:sink0_ready -> cmd_xbar_demux:src8_ready
	signal cmd_xbar_demux_src9_endofpacket                                                                        : std_logic;                      -- cmd_xbar_demux:src9_endofpacket -> cmd_xbar_mux_009:sink0_endofpacket
	signal cmd_xbar_demux_src9_valid                                                                              : std_logic;                      -- cmd_xbar_demux:src9_valid -> cmd_xbar_mux_009:sink0_valid
	signal cmd_xbar_demux_src9_startofpacket                                                                      : std_logic;                      -- cmd_xbar_demux:src9_startofpacket -> cmd_xbar_mux_009:sink0_startofpacket
	signal cmd_xbar_demux_src9_data                                                                               : std_logic_vector(99 downto 0);  -- cmd_xbar_demux:src9_data -> cmd_xbar_mux_009:sink0_data
	signal cmd_xbar_demux_src9_channel                                                                            : std_logic_vector(13 downto 0);  -- cmd_xbar_demux:src9_channel -> cmd_xbar_mux_009:sink0_channel
	signal cmd_xbar_demux_src9_ready                                                                              : std_logic;                      -- cmd_xbar_mux_009:sink0_ready -> cmd_xbar_demux:src9_ready
	signal cmd_xbar_demux_src10_endofpacket                                                                       : std_logic;                      -- cmd_xbar_demux:src10_endofpacket -> cmd_xbar_mux_010:sink0_endofpacket
	signal cmd_xbar_demux_src10_valid                                                                             : std_logic;                      -- cmd_xbar_demux:src10_valid -> cmd_xbar_mux_010:sink0_valid
	signal cmd_xbar_demux_src10_startofpacket                                                                     : std_logic;                      -- cmd_xbar_demux:src10_startofpacket -> cmd_xbar_mux_010:sink0_startofpacket
	signal cmd_xbar_demux_src10_data                                                                              : std_logic_vector(99 downto 0);  -- cmd_xbar_demux:src10_data -> cmd_xbar_mux_010:sink0_data
	signal cmd_xbar_demux_src10_channel                                                                           : std_logic_vector(13 downto 0);  -- cmd_xbar_demux:src10_channel -> cmd_xbar_mux_010:sink0_channel
	signal cmd_xbar_demux_src10_ready                                                                             : std_logic;                      -- cmd_xbar_mux_010:sink0_ready -> cmd_xbar_demux:src10_ready
	signal cmd_xbar_demux_src11_endofpacket                                                                       : std_logic;                      -- cmd_xbar_demux:src11_endofpacket -> cmd_xbar_mux_011:sink0_endofpacket
	signal cmd_xbar_demux_src11_valid                                                                             : std_logic;                      -- cmd_xbar_demux:src11_valid -> cmd_xbar_mux_011:sink0_valid
	signal cmd_xbar_demux_src11_startofpacket                                                                     : std_logic;                      -- cmd_xbar_demux:src11_startofpacket -> cmd_xbar_mux_011:sink0_startofpacket
	signal cmd_xbar_demux_src11_data                                                                              : std_logic_vector(99 downto 0);  -- cmd_xbar_demux:src11_data -> cmd_xbar_mux_011:sink0_data
	signal cmd_xbar_demux_src11_channel                                                                           : std_logic_vector(13 downto 0);  -- cmd_xbar_demux:src11_channel -> cmd_xbar_mux_011:sink0_channel
	signal cmd_xbar_demux_src11_ready                                                                             : std_logic;                      -- cmd_xbar_mux_011:sink0_ready -> cmd_xbar_demux:src11_ready
	signal cmd_xbar_demux_src12_endofpacket                                                                       : std_logic;                      -- cmd_xbar_demux:src12_endofpacket -> cmd_xbar_mux_012:sink0_endofpacket
	signal cmd_xbar_demux_src12_valid                                                                             : std_logic;                      -- cmd_xbar_demux:src12_valid -> cmd_xbar_mux_012:sink0_valid
	signal cmd_xbar_demux_src12_startofpacket                                                                     : std_logic;                      -- cmd_xbar_demux:src12_startofpacket -> cmd_xbar_mux_012:sink0_startofpacket
	signal cmd_xbar_demux_src12_data                                                                              : std_logic_vector(99 downto 0);  -- cmd_xbar_demux:src12_data -> cmd_xbar_mux_012:sink0_data
	signal cmd_xbar_demux_src12_channel                                                                           : std_logic_vector(13 downto 0);  -- cmd_xbar_demux:src12_channel -> cmd_xbar_mux_012:sink0_channel
	signal cmd_xbar_demux_src12_ready                                                                             : std_logic;                      -- cmd_xbar_mux_012:sink0_ready -> cmd_xbar_demux:src12_ready
	signal cmd_xbar_demux_src13_endofpacket                                                                       : std_logic;                      -- cmd_xbar_demux:src13_endofpacket -> cmd_xbar_mux_013:sink0_endofpacket
	signal cmd_xbar_demux_src13_valid                                                                             : std_logic;                      -- cmd_xbar_demux:src13_valid -> cmd_xbar_mux_013:sink0_valid
	signal cmd_xbar_demux_src13_startofpacket                                                                     : std_logic;                      -- cmd_xbar_demux:src13_startofpacket -> cmd_xbar_mux_013:sink0_startofpacket
	signal cmd_xbar_demux_src13_data                                                                              : std_logic_vector(99 downto 0);  -- cmd_xbar_demux:src13_data -> cmd_xbar_mux_013:sink0_data
	signal cmd_xbar_demux_src13_channel                                                                           : std_logic_vector(13 downto 0);  -- cmd_xbar_demux:src13_channel -> cmd_xbar_mux_013:sink0_channel
	signal cmd_xbar_demux_src13_ready                                                                             : std_logic;                      -- cmd_xbar_mux_013:sink0_ready -> cmd_xbar_demux:src13_ready
	signal cmd_xbar_demux_001_src0_endofpacket                                                                    : std_logic;                      -- cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	signal cmd_xbar_demux_001_src0_valid                                                                          : std_logic;                      -- cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	signal cmd_xbar_demux_001_src0_startofpacket                                                                  : std_logic;                      -- cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	signal cmd_xbar_demux_001_src0_data                                                                           : std_logic_vector(99 downto 0);  -- cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	signal cmd_xbar_demux_001_src0_channel                                                                        : std_logic_vector(13 downto 0);  -- cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	signal cmd_xbar_demux_001_src0_ready                                                                          : std_logic;                      -- cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	signal cmd_xbar_demux_001_src1_endofpacket                                                                    : std_logic;                      -- cmd_xbar_demux_001:src1_endofpacket -> cmd_xbar_mux_001:sink1_endofpacket
	signal cmd_xbar_demux_001_src1_valid                                                                          : std_logic;                      -- cmd_xbar_demux_001:src1_valid -> cmd_xbar_mux_001:sink1_valid
	signal cmd_xbar_demux_001_src1_startofpacket                                                                  : std_logic;                      -- cmd_xbar_demux_001:src1_startofpacket -> cmd_xbar_mux_001:sink1_startofpacket
	signal cmd_xbar_demux_001_src1_data                                                                           : std_logic_vector(99 downto 0);  -- cmd_xbar_demux_001:src1_data -> cmd_xbar_mux_001:sink1_data
	signal cmd_xbar_demux_001_src1_channel                                                                        : std_logic_vector(13 downto 0);  -- cmd_xbar_demux_001:src1_channel -> cmd_xbar_mux_001:sink1_channel
	signal cmd_xbar_demux_001_src1_ready                                                                          : std_logic;                      -- cmd_xbar_mux_001:sink1_ready -> cmd_xbar_demux_001:src1_ready
	signal cmd_xbar_demux_001_src2_endofpacket                                                                    : std_logic;                      -- cmd_xbar_demux_001:src2_endofpacket -> cmd_xbar_mux_002:sink1_endofpacket
	signal cmd_xbar_demux_001_src2_valid                                                                          : std_logic;                      -- cmd_xbar_demux_001:src2_valid -> cmd_xbar_mux_002:sink1_valid
	signal cmd_xbar_demux_001_src2_startofpacket                                                                  : std_logic;                      -- cmd_xbar_demux_001:src2_startofpacket -> cmd_xbar_mux_002:sink1_startofpacket
	signal cmd_xbar_demux_001_src2_data                                                                           : std_logic_vector(99 downto 0);  -- cmd_xbar_demux_001:src2_data -> cmd_xbar_mux_002:sink1_data
	signal cmd_xbar_demux_001_src2_channel                                                                        : std_logic_vector(13 downto 0);  -- cmd_xbar_demux_001:src2_channel -> cmd_xbar_mux_002:sink1_channel
	signal cmd_xbar_demux_001_src2_ready                                                                          : std_logic;                      -- cmd_xbar_mux_002:sink1_ready -> cmd_xbar_demux_001:src2_ready
	signal cmd_xbar_demux_001_src3_endofpacket                                                                    : std_logic;                      -- cmd_xbar_demux_001:src3_endofpacket -> cmd_xbar_mux_003:sink1_endofpacket
	signal cmd_xbar_demux_001_src3_valid                                                                          : std_logic;                      -- cmd_xbar_demux_001:src3_valid -> cmd_xbar_mux_003:sink1_valid
	signal cmd_xbar_demux_001_src3_startofpacket                                                                  : std_logic;                      -- cmd_xbar_demux_001:src3_startofpacket -> cmd_xbar_mux_003:sink1_startofpacket
	signal cmd_xbar_demux_001_src3_data                                                                           : std_logic_vector(99 downto 0);  -- cmd_xbar_demux_001:src3_data -> cmd_xbar_mux_003:sink1_data
	signal cmd_xbar_demux_001_src3_channel                                                                        : std_logic_vector(13 downto 0);  -- cmd_xbar_demux_001:src3_channel -> cmd_xbar_mux_003:sink1_channel
	signal cmd_xbar_demux_001_src3_ready                                                                          : std_logic;                      -- cmd_xbar_mux_003:sink1_ready -> cmd_xbar_demux_001:src3_ready
	signal cmd_xbar_demux_001_src4_endofpacket                                                                    : std_logic;                      -- cmd_xbar_demux_001:src4_endofpacket -> cmd_xbar_mux_004:sink1_endofpacket
	signal cmd_xbar_demux_001_src4_valid                                                                          : std_logic;                      -- cmd_xbar_demux_001:src4_valid -> cmd_xbar_mux_004:sink1_valid
	signal cmd_xbar_demux_001_src4_startofpacket                                                                  : std_logic;                      -- cmd_xbar_demux_001:src4_startofpacket -> cmd_xbar_mux_004:sink1_startofpacket
	signal cmd_xbar_demux_001_src4_data                                                                           : std_logic_vector(99 downto 0);  -- cmd_xbar_demux_001:src4_data -> cmd_xbar_mux_004:sink1_data
	signal cmd_xbar_demux_001_src4_channel                                                                        : std_logic_vector(13 downto 0);  -- cmd_xbar_demux_001:src4_channel -> cmd_xbar_mux_004:sink1_channel
	signal cmd_xbar_demux_001_src4_ready                                                                          : std_logic;                      -- cmd_xbar_mux_004:sink1_ready -> cmd_xbar_demux_001:src4_ready
	signal cmd_xbar_demux_001_src5_endofpacket                                                                    : std_logic;                      -- cmd_xbar_demux_001:src5_endofpacket -> cmd_xbar_mux_005:sink1_endofpacket
	signal cmd_xbar_demux_001_src5_valid                                                                          : std_logic;                      -- cmd_xbar_demux_001:src5_valid -> cmd_xbar_mux_005:sink1_valid
	signal cmd_xbar_demux_001_src5_startofpacket                                                                  : std_logic;                      -- cmd_xbar_demux_001:src5_startofpacket -> cmd_xbar_mux_005:sink1_startofpacket
	signal cmd_xbar_demux_001_src5_data                                                                           : std_logic_vector(99 downto 0);  -- cmd_xbar_demux_001:src5_data -> cmd_xbar_mux_005:sink1_data
	signal cmd_xbar_demux_001_src5_channel                                                                        : std_logic_vector(13 downto 0);  -- cmd_xbar_demux_001:src5_channel -> cmd_xbar_mux_005:sink1_channel
	signal cmd_xbar_demux_001_src5_ready                                                                          : std_logic;                      -- cmd_xbar_mux_005:sink1_ready -> cmd_xbar_demux_001:src5_ready
	signal cmd_xbar_demux_001_src6_endofpacket                                                                    : std_logic;                      -- cmd_xbar_demux_001:src6_endofpacket -> cmd_xbar_mux_006:sink1_endofpacket
	signal cmd_xbar_demux_001_src6_valid                                                                          : std_logic;                      -- cmd_xbar_demux_001:src6_valid -> cmd_xbar_mux_006:sink1_valid
	signal cmd_xbar_demux_001_src6_startofpacket                                                                  : std_logic;                      -- cmd_xbar_demux_001:src6_startofpacket -> cmd_xbar_mux_006:sink1_startofpacket
	signal cmd_xbar_demux_001_src6_data                                                                           : std_logic_vector(99 downto 0);  -- cmd_xbar_demux_001:src6_data -> cmd_xbar_mux_006:sink1_data
	signal cmd_xbar_demux_001_src6_channel                                                                        : std_logic_vector(13 downto 0);  -- cmd_xbar_demux_001:src6_channel -> cmd_xbar_mux_006:sink1_channel
	signal cmd_xbar_demux_001_src6_ready                                                                          : std_logic;                      -- cmd_xbar_mux_006:sink1_ready -> cmd_xbar_demux_001:src6_ready
	signal cmd_xbar_demux_001_src7_endofpacket                                                                    : std_logic;                      -- cmd_xbar_demux_001:src7_endofpacket -> cmd_xbar_mux_007:sink1_endofpacket
	signal cmd_xbar_demux_001_src7_valid                                                                          : std_logic;                      -- cmd_xbar_demux_001:src7_valid -> cmd_xbar_mux_007:sink1_valid
	signal cmd_xbar_demux_001_src7_startofpacket                                                                  : std_logic;                      -- cmd_xbar_demux_001:src7_startofpacket -> cmd_xbar_mux_007:sink1_startofpacket
	signal cmd_xbar_demux_001_src7_data                                                                           : std_logic_vector(99 downto 0);  -- cmd_xbar_demux_001:src7_data -> cmd_xbar_mux_007:sink1_data
	signal cmd_xbar_demux_001_src7_channel                                                                        : std_logic_vector(13 downto 0);  -- cmd_xbar_demux_001:src7_channel -> cmd_xbar_mux_007:sink1_channel
	signal cmd_xbar_demux_001_src7_ready                                                                          : std_logic;                      -- cmd_xbar_mux_007:sink1_ready -> cmd_xbar_demux_001:src7_ready
	signal cmd_xbar_demux_001_src8_endofpacket                                                                    : std_logic;                      -- cmd_xbar_demux_001:src8_endofpacket -> cmd_xbar_mux_008:sink1_endofpacket
	signal cmd_xbar_demux_001_src8_valid                                                                          : std_logic;                      -- cmd_xbar_demux_001:src8_valid -> cmd_xbar_mux_008:sink1_valid
	signal cmd_xbar_demux_001_src8_startofpacket                                                                  : std_logic;                      -- cmd_xbar_demux_001:src8_startofpacket -> cmd_xbar_mux_008:sink1_startofpacket
	signal cmd_xbar_demux_001_src8_data                                                                           : std_logic_vector(99 downto 0);  -- cmd_xbar_demux_001:src8_data -> cmd_xbar_mux_008:sink1_data
	signal cmd_xbar_demux_001_src8_channel                                                                        : std_logic_vector(13 downto 0);  -- cmd_xbar_demux_001:src8_channel -> cmd_xbar_mux_008:sink1_channel
	signal cmd_xbar_demux_001_src8_ready                                                                          : std_logic;                      -- cmd_xbar_mux_008:sink1_ready -> cmd_xbar_demux_001:src8_ready
	signal cmd_xbar_demux_001_src9_endofpacket                                                                    : std_logic;                      -- cmd_xbar_demux_001:src9_endofpacket -> cmd_xbar_mux_009:sink1_endofpacket
	signal cmd_xbar_demux_001_src9_valid                                                                          : std_logic;                      -- cmd_xbar_demux_001:src9_valid -> cmd_xbar_mux_009:sink1_valid
	signal cmd_xbar_demux_001_src9_startofpacket                                                                  : std_logic;                      -- cmd_xbar_demux_001:src9_startofpacket -> cmd_xbar_mux_009:sink1_startofpacket
	signal cmd_xbar_demux_001_src9_data                                                                           : std_logic_vector(99 downto 0);  -- cmd_xbar_demux_001:src9_data -> cmd_xbar_mux_009:sink1_data
	signal cmd_xbar_demux_001_src9_channel                                                                        : std_logic_vector(13 downto 0);  -- cmd_xbar_demux_001:src9_channel -> cmd_xbar_mux_009:sink1_channel
	signal cmd_xbar_demux_001_src9_ready                                                                          : std_logic;                      -- cmd_xbar_mux_009:sink1_ready -> cmd_xbar_demux_001:src9_ready
	signal cmd_xbar_demux_001_src10_endofpacket                                                                   : std_logic;                      -- cmd_xbar_demux_001:src10_endofpacket -> cmd_xbar_mux_010:sink1_endofpacket
	signal cmd_xbar_demux_001_src10_valid                                                                         : std_logic;                      -- cmd_xbar_demux_001:src10_valid -> cmd_xbar_mux_010:sink1_valid
	signal cmd_xbar_demux_001_src10_startofpacket                                                                 : std_logic;                      -- cmd_xbar_demux_001:src10_startofpacket -> cmd_xbar_mux_010:sink1_startofpacket
	signal cmd_xbar_demux_001_src10_data                                                                          : std_logic_vector(99 downto 0);  -- cmd_xbar_demux_001:src10_data -> cmd_xbar_mux_010:sink1_data
	signal cmd_xbar_demux_001_src10_channel                                                                       : std_logic_vector(13 downto 0);  -- cmd_xbar_demux_001:src10_channel -> cmd_xbar_mux_010:sink1_channel
	signal cmd_xbar_demux_001_src10_ready                                                                         : std_logic;                      -- cmd_xbar_mux_010:sink1_ready -> cmd_xbar_demux_001:src10_ready
	signal cmd_xbar_demux_001_src11_endofpacket                                                                   : std_logic;                      -- cmd_xbar_demux_001:src11_endofpacket -> cmd_xbar_mux_011:sink1_endofpacket
	signal cmd_xbar_demux_001_src11_valid                                                                         : std_logic;                      -- cmd_xbar_demux_001:src11_valid -> cmd_xbar_mux_011:sink1_valid
	signal cmd_xbar_demux_001_src11_startofpacket                                                                 : std_logic;                      -- cmd_xbar_demux_001:src11_startofpacket -> cmd_xbar_mux_011:sink1_startofpacket
	signal cmd_xbar_demux_001_src11_data                                                                          : std_logic_vector(99 downto 0);  -- cmd_xbar_demux_001:src11_data -> cmd_xbar_mux_011:sink1_data
	signal cmd_xbar_demux_001_src11_channel                                                                       : std_logic_vector(13 downto 0);  -- cmd_xbar_demux_001:src11_channel -> cmd_xbar_mux_011:sink1_channel
	signal cmd_xbar_demux_001_src11_ready                                                                         : std_logic;                      -- cmd_xbar_mux_011:sink1_ready -> cmd_xbar_demux_001:src11_ready
	signal cmd_xbar_demux_001_src12_endofpacket                                                                   : std_logic;                      -- cmd_xbar_demux_001:src12_endofpacket -> cmd_xbar_mux_012:sink1_endofpacket
	signal cmd_xbar_demux_001_src12_valid                                                                         : std_logic;                      -- cmd_xbar_demux_001:src12_valid -> cmd_xbar_mux_012:sink1_valid
	signal cmd_xbar_demux_001_src12_startofpacket                                                                 : std_logic;                      -- cmd_xbar_demux_001:src12_startofpacket -> cmd_xbar_mux_012:sink1_startofpacket
	signal cmd_xbar_demux_001_src12_data                                                                          : std_logic_vector(99 downto 0);  -- cmd_xbar_demux_001:src12_data -> cmd_xbar_mux_012:sink1_data
	signal cmd_xbar_demux_001_src12_channel                                                                       : std_logic_vector(13 downto 0);  -- cmd_xbar_demux_001:src12_channel -> cmd_xbar_mux_012:sink1_channel
	signal cmd_xbar_demux_001_src12_ready                                                                         : std_logic;                      -- cmd_xbar_mux_012:sink1_ready -> cmd_xbar_demux_001:src12_ready
	signal cmd_xbar_demux_001_src13_endofpacket                                                                   : std_logic;                      -- cmd_xbar_demux_001:src13_endofpacket -> cmd_xbar_mux_013:sink1_endofpacket
	signal cmd_xbar_demux_001_src13_valid                                                                         : std_logic;                      -- cmd_xbar_demux_001:src13_valid -> cmd_xbar_mux_013:sink1_valid
	signal cmd_xbar_demux_001_src13_startofpacket                                                                 : std_logic;                      -- cmd_xbar_demux_001:src13_startofpacket -> cmd_xbar_mux_013:sink1_startofpacket
	signal cmd_xbar_demux_001_src13_data                                                                          : std_logic_vector(99 downto 0);  -- cmd_xbar_demux_001:src13_data -> cmd_xbar_mux_013:sink1_data
	signal cmd_xbar_demux_001_src13_channel                                                                       : std_logic_vector(13 downto 0);  -- cmd_xbar_demux_001:src13_channel -> cmd_xbar_mux_013:sink1_channel
	signal cmd_xbar_demux_001_src13_ready                                                                         : std_logic;                      -- cmd_xbar_mux_013:sink1_ready -> cmd_xbar_demux_001:src13_ready
	signal rsp_xbar_demux_src0_endofpacket                                                                        : std_logic;                      -- rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	signal rsp_xbar_demux_src0_valid                                                                              : std_logic;                      -- rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	signal rsp_xbar_demux_src0_startofpacket                                                                      : std_logic;                      -- rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	signal rsp_xbar_demux_src0_data                                                                               : std_logic_vector(99 downto 0);  -- rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	signal rsp_xbar_demux_src0_channel                                                                            : std_logic_vector(13 downto 0);  -- rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	signal rsp_xbar_demux_src0_ready                                                                              : std_logic;                      -- rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	signal rsp_xbar_demux_src1_endofpacket                                                                        : std_logic;                      -- rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	signal rsp_xbar_demux_src1_valid                                                                              : std_logic;                      -- rsp_xbar_demux:src1_valid -> rsp_xbar_mux_001:sink0_valid
	signal rsp_xbar_demux_src1_startofpacket                                                                      : std_logic;                      -- rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	signal rsp_xbar_demux_src1_data                                                                               : std_logic_vector(99 downto 0);  -- rsp_xbar_demux:src1_data -> rsp_xbar_mux_001:sink0_data
	signal rsp_xbar_demux_src1_channel                                                                            : std_logic_vector(13 downto 0);  -- rsp_xbar_demux:src1_channel -> rsp_xbar_mux_001:sink0_channel
	signal rsp_xbar_demux_src1_ready                                                                              : std_logic;                      -- rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux:src1_ready
	signal rsp_xbar_demux_001_src0_endofpacket                                                                    : std_logic;                      -- rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	signal rsp_xbar_demux_001_src0_valid                                                                          : std_logic;                      -- rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	signal rsp_xbar_demux_001_src0_startofpacket                                                                  : std_logic;                      -- rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	signal rsp_xbar_demux_001_src0_data                                                                           : std_logic_vector(99 downto 0);  -- rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	signal rsp_xbar_demux_001_src0_channel                                                                        : std_logic_vector(13 downto 0);  -- rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	signal rsp_xbar_demux_001_src0_ready                                                                          : std_logic;                      -- rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	signal rsp_xbar_demux_001_src1_endofpacket                                                                    : std_logic;                      -- rsp_xbar_demux_001:src1_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	signal rsp_xbar_demux_001_src1_valid                                                                          : std_logic;                      -- rsp_xbar_demux_001:src1_valid -> rsp_xbar_mux_001:sink1_valid
	signal rsp_xbar_demux_001_src1_startofpacket                                                                  : std_logic;                      -- rsp_xbar_demux_001:src1_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	signal rsp_xbar_demux_001_src1_data                                                                           : std_logic_vector(99 downto 0);  -- rsp_xbar_demux_001:src1_data -> rsp_xbar_mux_001:sink1_data
	signal rsp_xbar_demux_001_src1_channel                                                                        : std_logic_vector(13 downto 0);  -- rsp_xbar_demux_001:src1_channel -> rsp_xbar_mux_001:sink1_channel
	signal rsp_xbar_demux_001_src1_ready                                                                          : std_logic;                      -- rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_001:src1_ready
	signal rsp_xbar_demux_002_src0_endofpacket                                                                    : std_logic;                      -- rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux:sink2_endofpacket
	signal rsp_xbar_demux_002_src0_valid                                                                          : std_logic;                      -- rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux:sink2_valid
	signal rsp_xbar_demux_002_src0_startofpacket                                                                  : std_logic;                      -- rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux:sink2_startofpacket
	signal rsp_xbar_demux_002_src0_data                                                                           : std_logic_vector(99 downto 0);  -- rsp_xbar_demux_002:src0_data -> rsp_xbar_mux:sink2_data
	signal rsp_xbar_demux_002_src0_channel                                                                        : std_logic_vector(13 downto 0);  -- rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux:sink2_channel
	signal rsp_xbar_demux_002_src0_ready                                                                          : std_logic;                      -- rsp_xbar_mux:sink2_ready -> rsp_xbar_demux_002:src0_ready
	signal rsp_xbar_demux_002_src1_endofpacket                                                                    : std_logic;                      -- rsp_xbar_demux_002:src1_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	signal rsp_xbar_demux_002_src1_valid                                                                          : std_logic;                      -- rsp_xbar_demux_002:src1_valid -> rsp_xbar_mux_001:sink2_valid
	signal rsp_xbar_demux_002_src1_startofpacket                                                                  : std_logic;                      -- rsp_xbar_demux_002:src1_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	signal rsp_xbar_demux_002_src1_data                                                                           : std_logic_vector(99 downto 0);  -- rsp_xbar_demux_002:src1_data -> rsp_xbar_mux_001:sink2_data
	signal rsp_xbar_demux_002_src1_channel                                                                        : std_logic_vector(13 downto 0);  -- rsp_xbar_demux_002:src1_channel -> rsp_xbar_mux_001:sink2_channel
	signal rsp_xbar_demux_002_src1_ready                                                                          : std_logic;                      -- rsp_xbar_mux_001:sink2_ready -> rsp_xbar_demux_002:src1_ready
	signal rsp_xbar_demux_003_src0_endofpacket                                                                    : std_logic;                      -- rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux:sink3_endofpacket
	signal rsp_xbar_demux_003_src0_valid                                                                          : std_logic;                      -- rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux:sink3_valid
	signal rsp_xbar_demux_003_src0_startofpacket                                                                  : std_logic;                      -- rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux:sink3_startofpacket
	signal rsp_xbar_demux_003_src0_data                                                                           : std_logic_vector(99 downto 0);  -- rsp_xbar_demux_003:src0_data -> rsp_xbar_mux:sink3_data
	signal rsp_xbar_demux_003_src0_channel                                                                        : std_logic_vector(13 downto 0);  -- rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux:sink3_channel
	signal rsp_xbar_demux_003_src0_ready                                                                          : std_logic;                      -- rsp_xbar_mux:sink3_ready -> rsp_xbar_demux_003:src0_ready
	signal rsp_xbar_demux_003_src1_endofpacket                                                                    : std_logic;                      -- rsp_xbar_demux_003:src1_endofpacket -> rsp_xbar_mux_001:sink3_endofpacket
	signal rsp_xbar_demux_003_src1_valid                                                                          : std_logic;                      -- rsp_xbar_demux_003:src1_valid -> rsp_xbar_mux_001:sink3_valid
	signal rsp_xbar_demux_003_src1_startofpacket                                                                  : std_logic;                      -- rsp_xbar_demux_003:src1_startofpacket -> rsp_xbar_mux_001:sink3_startofpacket
	signal rsp_xbar_demux_003_src1_data                                                                           : std_logic_vector(99 downto 0);  -- rsp_xbar_demux_003:src1_data -> rsp_xbar_mux_001:sink3_data
	signal rsp_xbar_demux_003_src1_channel                                                                        : std_logic_vector(13 downto 0);  -- rsp_xbar_demux_003:src1_channel -> rsp_xbar_mux_001:sink3_channel
	signal rsp_xbar_demux_003_src1_ready                                                                          : std_logic;                      -- rsp_xbar_mux_001:sink3_ready -> rsp_xbar_demux_003:src1_ready
	signal rsp_xbar_demux_004_src0_endofpacket                                                                    : std_logic;                      -- rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux:sink4_endofpacket
	signal rsp_xbar_demux_004_src0_valid                                                                          : std_logic;                      -- rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux:sink4_valid
	signal rsp_xbar_demux_004_src0_startofpacket                                                                  : std_logic;                      -- rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux:sink4_startofpacket
	signal rsp_xbar_demux_004_src0_data                                                                           : std_logic_vector(99 downto 0);  -- rsp_xbar_demux_004:src0_data -> rsp_xbar_mux:sink4_data
	signal rsp_xbar_demux_004_src0_channel                                                                        : std_logic_vector(13 downto 0);  -- rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux:sink4_channel
	signal rsp_xbar_demux_004_src0_ready                                                                          : std_logic;                      -- rsp_xbar_mux:sink4_ready -> rsp_xbar_demux_004:src0_ready
	signal rsp_xbar_demux_004_src1_endofpacket                                                                    : std_logic;                      -- rsp_xbar_demux_004:src1_endofpacket -> rsp_xbar_mux_001:sink4_endofpacket
	signal rsp_xbar_demux_004_src1_valid                                                                          : std_logic;                      -- rsp_xbar_demux_004:src1_valid -> rsp_xbar_mux_001:sink4_valid
	signal rsp_xbar_demux_004_src1_startofpacket                                                                  : std_logic;                      -- rsp_xbar_demux_004:src1_startofpacket -> rsp_xbar_mux_001:sink4_startofpacket
	signal rsp_xbar_demux_004_src1_data                                                                           : std_logic_vector(99 downto 0);  -- rsp_xbar_demux_004:src1_data -> rsp_xbar_mux_001:sink4_data
	signal rsp_xbar_demux_004_src1_channel                                                                        : std_logic_vector(13 downto 0);  -- rsp_xbar_demux_004:src1_channel -> rsp_xbar_mux_001:sink4_channel
	signal rsp_xbar_demux_004_src1_ready                                                                          : std_logic;                      -- rsp_xbar_mux_001:sink4_ready -> rsp_xbar_demux_004:src1_ready
	signal rsp_xbar_demux_005_src0_endofpacket                                                                    : std_logic;                      -- rsp_xbar_demux_005:src0_endofpacket -> rsp_xbar_mux:sink5_endofpacket
	signal rsp_xbar_demux_005_src0_valid                                                                          : std_logic;                      -- rsp_xbar_demux_005:src0_valid -> rsp_xbar_mux:sink5_valid
	signal rsp_xbar_demux_005_src0_startofpacket                                                                  : std_logic;                      -- rsp_xbar_demux_005:src0_startofpacket -> rsp_xbar_mux:sink5_startofpacket
	signal rsp_xbar_demux_005_src0_data                                                                           : std_logic_vector(99 downto 0);  -- rsp_xbar_demux_005:src0_data -> rsp_xbar_mux:sink5_data
	signal rsp_xbar_demux_005_src0_channel                                                                        : std_logic_vector(13 downto 0);  -- rsp_xbar_demux_005:src0_channel -> rsp_xbar_mux:sink5_channel
	signal rsp_xbar_demux_005_src0_ready                                                                          : std_logic;                      -- rsp_xbar_mux:sink5_ready -> rsp_xbar_demux_005:src0_ready
	signal rsp_xbar_demux_005_src1_endofpacket                                                                    : std_logic;                      -- rsp_xbar_demux_005:src1_endofpacket -> rsp_xbar_mux_001:sink5_endofpacket
	signal rsp_xbar_demux_005_src1_valid                                                                          : std_logic;                      -- rsp_xbar_demux_005:src1_valid -> rsp_xbar_mux_001:sink5_valid
	signal rsp_xbar_demux_005_src1_startofpacket                                                                  : std_logic;                      -- rsp_xbar_demux_005:src1_startofpacket -> rsp_xbar_mux_001:sink5_startofpacket
	signal rsp_xbar_demux_005_src1_data                                                                           : std_logic_vector(99 downto 0);  -- rsp_xbar_demux_005:src1_data -> rsp_xbar_mux_001:sink5_data
	signal rsp_xbar_demux_005_src1_channel                                                                        : std_logic_vector(13 downto 0);  -- rsp_xbar_demux_005:src1_channel -> rsp_xbar_mux_001:sink5_channel
	signal rsp_xbar_demux_005_src1_ready                                                                          : std_logic;                      -- rsp_xbar_mux_001:sink5_ready -> rsp_xbar_demux_005:src1_ready
	signal rsp_xbar_demux_006_src0_endofpacket                                                                    : std_logic;                      -- rsp_xbar_demux_006:src0_endofpacket -> rsp_xbar_mux:sink6_endofpacket
	signal rsp_xbar_demux_006_src0_valid                                                                          : std_logic;                      -- rsp_xbar_demux_006:src0_valid -> rsp_xbar_mux:sink6_valid
	signal rsp_xbar_demux_006_src0_startofpacket                                                                  : std_logic;                      -- rsp_xbar_demux_006:src0_startofpacket -> rsp_xbar_mux:sink6_startofpacket
	signal rsp_xbar_demux_006_src0_data                                                                           : std_logic_vector(99 downto 0);  -- rsp_xbar_demux_006:src0_data -> rsp_xbar_mux:sink6_data
	signal rsp_xbar_demux_006_src0_channel                                                                        : std_logic_vector(13 downto 0);  -- rsp_xbar_demux_006:src0_channel -> rsp_xbar_mux:sink6_channel
	signal rsp_xbar_demux_006_src0_ready                                                                          : std_logic;                      -- rsp_xbar_mux:sink6_ready -> rsp_xbar_demux_006:src0_ready
	signal rsp_xbar_demux_006_src1_endofpacket                                                                    : std_logic;                      -- rsp_xbar_demux_006:src1_endofpacket -> rsp_xbar_mux_001:sink6_endofpacket
	signal rsp_xbar_demux_006_src1_valid                                                                          : std_logic;                      -- rsp_xbar_demux_006:src1_valid -> rsp_xbar_mux_001:sink6_valid
	signal rsp_xbar_demux_006_src1_startofpacket                                                                  : std_logic;                      -- rsp_xbar_demux_006:src1_startofpacket -> rsp_xbar_mux_001:sink6_startofpacket
	signal rsp_xbar_demux_006_src1_data                                                                           : std_logic_vector(99 downto 0);  -- rsp_xbar_demux_006:src1_data -> rsp_xbar_mux_001:sink6_data
	signal rsp_xbar_demux_006_src1_channel                                                                        : std_logic_vector(13 downto 0);  -- rsp_xbar_demux_006:src1_channel -> rsp_xbar_mux_001:sink6_channel
	signal rsp_xbar_demux_006_src1_ready                                                                          : std_logic;                      -- rsp_xbar_mux_001:sink6_ready -> rsp_xbar_demux_006:src1_ready
	signal rsp_xbar_demux_007_src0_endofpacket                                                                    : std_logic;                      -- rsp_xbar_demux_007:src0_endofpacket -> rsp_xbar_mux:sink7_endofpacket
	signal rsp_xbar_demux_007_src0_valid                                                                          : std_logic;                      -- rsp_xbar_demux_007:src0_valid -> rsp_xbar_mux:sink7_valid
	signal rsp_xbar_demux_007_src0_startofpacket                                                                  : std_logic;                      -- rsp_xbar_demux_007:src0_startofpacket -> rsp_xbar_mux:sink7_startofpacket
	signal rsp_xbar_demux_007_src0_data                                                                           : std_logic_vector(99 downto 0);  -- rsp_xbar_demux_007:src0_data -> rsp_xbar_mux:sink7_data
	signal rsp_xbar_demux_007_src0_channel                                                                        : std_logic_vector(13 downto 0);  -- rsp_xbar_demux_007:src0_channel -> rsp_xbar_mux:sink7_channel
	signal rsp_xbar_demux_007_src0_ready                                                                          : std_logic;                      -- rsp_xbar_mux:sink7_ready -> rsp_xbar_demux_007:src0_ready
	signal rsp_xbar_demux_007_src1_endofpacket                                                                    : std_logic;                      -- rsp_xbar_demux_007:src1_endofpacket -> rsp_xbar_mux_001:sink7_endofpacket
	signal rsp_xbar_demux_007_src1_valid                                                                          : std_logic;                      -- rsp_xbar_demux_007:src1_valid -> rsp_xbar_mux_001:sink7_valid
	signal rsp_xbar_demux_007_src1_startofpacket                                                                  : std_logic;                      -- rsp_xbar_demux_007:src1_startofpacket -> rsp_xbar_mux_001:sink7_startofpacket
	signal rsp_xbar_demux_007_src1_data                                                                           : std_logic_vector(99 downto 0);  -- rsp_xbar_demux_007:src1_data -> rsp_xbar_mux_001:sink7_data
	signal rsp_xbar_demux_007_src1_channel                                                                        : std_logic_vector(13 downto 0);  -- rsp_xbar_demux_007:src1_channel -> rsp_xbar_mux_001:sink7_channel
	signal rsp_xbar_demux_007_src1_ready                                                                          : std_logic;                      -- rsp_xbar_mux_001:sink7_ready -> rsp_xbar_demux_007:src1_ready
	signal rsp_xbar_demux_008_src0_endofpacket                                                                    : std_logic;                      -- rsp_xbar_demux_008:src0_endofpacket -> rsp_xbar_mux:sink8_endofpacket
	signal rsp_xbar_demux_008_src0_valid                                                                          : std_logic;                      -- rsp_xbar_demux_008:src0_valid -> rsp_xbar_mux:sink8_valid
	signal rsp_xbar_demux_008_src0_startofpacket                                                                  : std_logic;                      -- rsp_xbar_demux_008:src0_startofpacket -> rsp_xbar_mux:sink8_startofpacket
	signal rsp_xbar_demux_008_src0_data                                                                           : std_logic_vector(99 downto 0);  -- rsp_xbar_demux_008:src0_data -> rsp_xbar_mux:sink8_data
	signal rsp_xbar_demux_008_src0_channel                                                                        : std_logic_vector(13 downto 0);  -- rsp_xbar_demux_008:src0_channel -> rsp_xbar_mux:sink8_channel
	signal rsp_xbar_demux_008_src0_ready                                                                          : std_logic;                      -- rsp_xbar_mux:sink8_ready -> rsp_xbar_demux_008:src0_ready
	signal rsp_xbar_demux_008_src1_endofpacket                                                                    : std_logic;                      -- rsp_xbar_demux_008:src1_endofpacket -> rsp_xbar_mux_001:sink8_endofpacket
	signal rsp_xbar_demux_008_src1_valid                                                                          : std_logic;                      -- rsp_xbar_demux_008:src1_valid -> rsp_xbar_mux_001:sink8_valid
	signal rsp_xbar_demux_008_src1_startofpacket                                                                  : std_logic;                      -- rsp_xbar_demux_008:src1_startofpacket -> rsp_xbar_mux_001:sink8_startofpacket
	signal rsp_xbar_demux_008_src1_data                                                                           : std_logic_vector(99 downto 0);  -- rsp_xbar_demux_008:src1_data -> rsp_xbar_mux_001:sink8_data
	signal rsp_xbar_demux_008_src1_channel                                                                        : std_logic_vector(13 downto 0);  -- rsp_xbar_demux_008:src1_channel -> rsp_xbar_mux_001:sink8_channel
	signal rsp_xbar_demux_008_src1_ready                                                                          : std_logic;                      -- rsp_xbar_mux_001:sink8_ready -> rsp_xbar_demux_008:src1_ready
	signal rsp_xbar_demux_009_src0_endofpacket                                                                    : std_logic;                      -- rsp_xbar_demux_009:src0_endofpacket -> rsp_xbar_mux:sink9_endofpacket
	signal rsp_xbar_demux_009_src0_valid                                                                          : std_logic;                      -- rsp_xbar_demux_009:src0_valid -> rsp_xbar_mux:sink9_valid
	signal rsp_xbar_demux_009_src0_startofpacket                                                                  : std_logic;                      -- rsp_xbar_demux_009:src0_startofpacket -> rsp_xbar_mux:sink9_startofpacket
	signal rsp_xbar_demux_009_src0_data                                                                           : std_logic_vector(99 downto 0);  -- rsp_xbar_demux_009:src0_data -> rsp_xbar_mux:sink9_data
	signal rsp_xbar_demux_009_src0_channel                                                                        : std_logic_vector(13 downto 0);  -- rsp_xbar_demux_009:src0_channel -> rsp_xbar_mux:sink9_channel
	signal rsp_xbar_demux_009_src0_ready                                                                          : std_logic;                      -- rsp_xbar_mux:sink9_ready -> rsp_xbar_demux_009:src0_ready
	signal rsp_xbar_demux_009_src1_endofpacket                                                                    : std_logic;                      -- rsp_xbar_demux_009:src1_endofpacket -> rsp_xbar_mux_001:sink9_endofpacket
	signal rsp_xbar_demux_009_src1_valid                                                                          : std_logic;                      -- rsp_xbar_demux_009:src1_valid -> rsp_xbar_mux_001:sink9_valid
	signal rsp_xbar_demux_009_src1_startofpacket                                                                  : std_logic;                      -- rsp_xbar_demux_009:src1_startofpacket -> rsp_xbar_mux_001:sink9_startofpacket
	signal rsp_xbar_demux_009_src1_data                                                                           : std_logic_vector(99 downto 0);  -- rsp_xbar_demux_009:src1_data -> rsp_xbar_mux_001:sink9_data
	signal rsp_xbar_demux_009_src1_channel                                                                        : std_logic_vector(13 downto 0);  -- rsp_xbar_demux_009:src1_channel -> rsp_xbar_mux_001:sink9_channel
	signal rsp_xbar_demux_009_src1_ready                                                                          : std_logic;                      -- rsp_xbar_mux_001:sink9_ready -> rsp_xbar_demux_009:src1_ready
	signal rsp_xbar_demux_010_src0_endofpacket                                                                    : std_logic;                      -- rsp_xbar_demux_010:src0_endofpacket -> rsp_xbar_mux:sink10_endofpacket
	signal rsp_xbar_demux_010_src0_valid                                                                          : std_logic;                      -- rsp_xbar_demux_010:src0_valid -> rsp_xbar_mux:sink10_valid
	signal rsp_xbar_demux_010_src0_startofpacket                                                                  : std_logic;                      -- rsp_xbar_demux_010:src0_startofpacket -> rsp_xbar_mux:sink10_startofpacket
	signal rsp_xbar_demux_010_src0_data                                                                           : std_logic_vector(99 downto 0);  -- rsp_xbar_demux_010:src0_data -> rsp_xbar_mux:sink10_data
	signal rsp_xbar_demux_010_src0_channel                                                                        : std_logic_vector(13 downto 0);  -- rsp_xbar_demux_010:src0_channel -> rsp_xbar_mux:sink10_channel
	signal rsp_xbar_demux_010_src0_ready                                                                          : std_logic;                      -- rsp_xbar_mux:sink10_ready -> rsp_xbar_demux_010:src0_ready
	signal rsp_xbar_demux_010_src1_endofpacket                                                                    : std_logic;                      -- rsp_xbar_demux_010:src1_endofpacket -> rsp_xbar_mux_001:sink10_endofpacket
	signal rsp_xbar_demux_010_src1_valid                                                                          : std_logic;                      -- rsp_xbar_demux_010:src1_valid -> rsp_xbar_mux_001:sink10_valid
	signal rsp_xbar_demux_010_src1_startofpacket                                                                  : std_logic;                      -- rsp_xbar_demux_010:src1_startofpacket -> rsp_xbar_mux_001:sink10_startofpacket
	signal rsp_xbar_demux_010_src1_data                                                                           : std_logic_vector(99 downto 0);  -- rsp_xbar_demux_010:src1_data -> rsp_xbar_mux_001:sink10_data
	signal rsp_xbar_demux_010_src1_channel                                                                        : std_logic_vector(13 downto 0);  -- rsp_xbar_demux_010:src1_channel -> rsp_xbar_mux_001:sink10_channel
	signal rsp_xbar_demux_010_src1_ready                                                                          : std_logic;                      -- rsp_xbar_mux_001:sink10_ready -> rsp_xbar_demux_010:src1_ready
	signal rsp_xbar_demux_011_src0_endofpacket                                                                    : std_logic;                      -- rsp_xbar_demux_011:src0_endofpacket -> rsp_xbar_mux:sink11_endofpacket
	signal rsp_xbar_demux_011_src0_valid                                                                          : std_logic;                      -- rsp_xbar_demux_011:src0_valid -> rsp_xbar_mux:sink11_valid
	signal rsp_xbar_demux_011_src0_startofpacket                                                                  : std_logic;                      -- rsp_xbar_demux_011:src0_startofpacket -> rsp_xbar_mux:sink11_startofpacket
	signal rsp_xbar_demux_011_src0_data                                                                           : std_logic_vector(99 downto 0);  -- rsp_xbar_demux_011:src0_data -> rsp_xbar_mux:sink11_data
	signal rsp_xbar_demux_011_src0_channel                                                                        : std_logic_vector(13 downto 0);  -- rsp_xbar_demux_011:src0_channel -> rsp_xbar_mux:sink11_channel
	signal rsp_xbar_demux_011_src0_ready                                                                          : std_logic;                      -- rsp_xbar_mux:sink11_ready -> rsp_xbar_demux_011:src0_ready
	signal rsp_xbar_demux_011_src1_endofpacket                                                                    : std_logic;                      -- rsp_xbar_demux_011:src1_endofpacket -> rsp_xbar_mux_001:sink11_endofpacket
	signal rsp_xbar_demux_011_src1_valid                                                                          : std_logic;                      -- rsp_xbar_demux_011:src1_valid -> rsp_xbar_mux_001:sink11_valid
	signal rsp_xbar_demux_011_src1_startofpacket                                                                  : std_logic;                      -- rsp_xbar_demux_011:src1_startofpacket -> rsp_xbar_mux_001:sink11_startofpacket
	signal rsp_xbar_demux_011_src1_data                                                                           : std_logic_vector(99 downto 0);  -- rsp_xbar_demux_011:src1_data -> rsp_xbar_mux_001:sink11_data
	signal rsp_xbar_demux_011_src1_channel                                                                        : std_logic_vector(13 downto 0);  -- rsp_xbar_demux_011:src1_channel -> rsp_xbar_mux_001:sink11_channel
	signal rsp_xbar_demux_011_src1_ready                                                                          : std_logic;                      -- rsp_xbar_mux_001:sink11_ready -> rsp_xbar_demux_011:src1_ready
	signal rsp_xbar_demux_012_src0_endofpacket                                                                    : std_logic;                      -- rsp_xbar_demux_012:src0_endofpacket -> rsp_xbar_mux:sink12_endofpacket
	signal rsp_xbar_demux_012_src0_valid                                                                          : std_logic;                      -- rsp_xbar_demux_012:src0_valid -> rsp_xbar_mux:sink12_valid
	signal rsp_xbar_demux_012_src0_startofpacket                                                                  : std_logic;                      -- rsp_xbar_demux_012:src0_startofpacket -> rsp_xbar_mux:sink12_startofpacket
	signal rsp_xbar_demux_012_src0_data                                                                           : std_logic_vector(99 downto 0);  -- rsp_xbar_demux_012:src0_data -> rsp_xbar_mux:sink12_data
	signal rsp_xbar_demux_012_src0_channel                                                                        : std_logic_vector(13 downto 0);  -- rsp_xbar_demux_012:src0_channel -> rsp_xbar_mux:sink12_channel
	signal rsp_xbar_demux_012_src0_ready                                                                          : std_logic;                      -- rsp_xbar_mux:sink12_ready -> rsp_xbar_demux_012:src0_ready
	signal rsp_xbar_demux_012_src1_endofpacket                                                                    : std_logic;                      -- rsp_xbar_demux_012:src1_endofpacket -> rsp_xbar_mux_001:sink12_endofpacket
	signal rsp_xbar_demux_012_src1_valid                                                                          : std_logic;                      -- rsp_xbar_demux_012:src1_valid -> rsp_xbar_mux_001:sink12_valid
	signal rsp_xbar_demux_012_src1_startofpacket                                                                  : std_logic;                      -- rsp_xbar_demux_012:src1_startofpacket -> rsp_xbar_mux_001:sink12_startofpacket
	signal rsp_xbar_demux_012_src1_data                                                                           : std_logic_vector(99 downto 0);  -- rsp_xbar_demux_012:src1_data -> rsp_xbar_mux_001:sink12_data
	signal rsp_xbar_demux_012_src1_channel                                                                        : std_logic_vector(13 downto 0);  -- rsp_xbar_demux_012:src1_channel -> rsp_xbar_mux_001:sink12_channel
	signal rsp_xbar_demux_012_src1_ready                                                                          : std_logic;                      -- rsp_xbar_mux_001:sink12_ready -> rsp_xbar_demux_012:src1_ready
	signal rsp_xbar_demux_013_src0_endofpacket                                                                    : std_logic;                      -- rsp_xbar_demux_013:src0_endofpacket -> rsp_xbar_mux:sink13_endofpacket
	signal rsp_xbar_demux_013_src0_valid                                                                          : std_logic;                      -- rsp_xbar_demux_013:src0_valid -> rsp_xbar_mux:sink13_valid
	signal rsp_xbar_demux_013_src0_startofpacket                                                                  : std_logic;                      -- rsp_xbar_demux_013:src0_startofpacket -> rsp_xbar_mux:sink13_startofpacket
	signal rsp_xbar_demux_013_src0_data                                                                           : std_logic_vector(99 downto 0);  -- rsp_xbar_demux_013:src0_data -> rsp_xbar_mux:sink13_data
	signal rsp_xbar_demux_013_src0_channel                                                                        : std_logic_vector(13 downto 0);  -- rsp_xbar_demux_013:src0_channel -> rsp_xbar_mux:sink13_channel
	signal rsp_xbar_demux_013_src0_ready                                                                          : std_logic;                      -- rsp_xbar_mux:sink13_ready -> rsp_xbar_demux_013:src0_ready
	signal rsp_xbar_demux_013_src1_endofpacket                                                                    : std_logic;                      -- rsp_xbar_demux_013:src1_endofpacket -> rsp_xbar_mux_001:sink13_endofpacket
	signal rsp_xbar_demux_013_src1_valid                                                                          : std_logic;                      -- rsp_xbar_demux_013:src1_valid -> rsp_xbar_mux_001:sink13_valid
	signal rsp_xbar_demux_013_src1_startofpacket                                                                  : std_logic;                      -- rsp_xbar_demux_013:src1_startofpacket -> rsp_xbar_mux_001:sink13_startofpacket
	signal rsp_xbar_demux_013_src1_data                                                                           : std_logic_vector(99 downto 0);  -- rsp_xbar_demux_013:src1_data -> rsp_xbar_mux_001:sink13_data
	signal rsp_xbar_demux_013_src1_channel                                                                        : std_logic_vector(13 downto 0);  -- rsp_xbar_demux_013:src1_channel -> rsp_xbar_mux_001:sink13_channel
	signal rsp_xbar_demux_013_src1_ready                                                                          : std_logic;                      -- rsp_xbar_mux_001:sink13_ready -> rsp_xbar_demux_013:src1_ready
	signal addr_router_src_endofpacket                                                                            : std_logic;                      -- addr_router:src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	signal addr_router_src_valid                                                                                  : std_logic;                      -- addr_router:src_valid -> cmd_xbar_demux:sink_valid
	signal addr_router_src_startofpacket                                                                          : std_logic;                      -- addr_router:src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	signal addr_router_src_data                                                                                   : std_logic_vector(99 downto 0);  -- addr_router:src_data -> cmd_xbar_demux:sink_data
	signal addr_router_src_channel                                                                                : std_logic_vector(13 downto 0);  -- addr_router:src_channel -> cmd_xbar_demux:sink_channel
	signal addr_router_src_ready                                                                                  : std_logic;                      -- cmd_xbar_demux:sink_ready -> addr_router:src_ready
	signal rsp_xbar_mux_src_endofpacket                                                                           : std_logic;                      -- rsp_xbar_mux:src_endofpacket -> nios2_qsys_grms_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	signal rsp_xbar_mux_src_valid                                                                                 : std_logic;                      -- rsp_xbar_mux:src_valid -> nios2_qsys_grms_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	signal rsp_xbar_mux_src_startofpacket                                                                         : std_logic;                      -- rsp_xbar_mux:src_startofpacket -> nios2_qsys_grms_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	signal rsp_xbar_mux_src_data                                                                                  : std_logic_vector(99 downto 0);  -- rsp_xbar_mux:src_data -> nios2_qsys_grms_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	signal rsp_xbar_mux_src_channel                                                                               : std_logic_vector(13 downto 0);  -- rsp_xbar_mux:src_channel -> nios2_qsys_grms_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	signal rsp_xbar_mux_src_ready                                                                                 : std_logic;                      -- nios2_qsys_grms_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux:src_ready
	signal addr_router_001_src_endofpacket                                                                        : std_logic;                      -- addr_router_001:src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	signal addr_router_001_src_valid                                                                              : std_logic;                      -- addr_router_001:src_valid -> cmd_xbar_demux_001:sink_valid
	signal addr_router_001_src_startofpacket                                                                      : std_logic;                      -- addr_router_001:src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	signal addr_router_001_src_data                                                                               : std_logic_vector(99 downto 0);  -- addr_router_001:src_data -> cmd_xbar_demux_001:sink_data
	signal addr_router_001_src_channel                                                                            : std_logic_vector(13 downto 0);  -- addr_router_001:src_channel -> cmd_xbar_demux_001:sink_channel
	signal addr_router_001_src_ready                                                                              : std_logic;                      -- cmd_xbar_demux_001:sink_ready -> addr_router_001:src_ready
	signal rsp_xbar_mux_001_src_endofpacket                                                                       : std_logic;                      -- rsp_xbar_mux_001:src_endofpacket -> nios2_qsys_grms_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	signal rsp_xbar_mux_001_src_valid                                                                             : std_logic;                      -- rsp_xbar_mux_001:src_valid -> nios2_qsys_grms_data_master_translator_avalon_universal_master_0_agent:rp_valid
	signal rsp_xbar_mux_001_src_startofpacket                                                                     : std_logic;                      -- rsp_xbar_mux_001:src_startofpacket -> nios2_qsys_grms_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	signal rsp_xbar_mux_001_src_data                                                                              : std_logic_vector(99 downto 0);  -- rsp_xbar_mux_001:src_data -> nios2_qsys_grms_data_master_translator_avalon_universal_master_0_agent:rp_data
	signal rsp_xbar_mux_001_src_channel                                                                           : std_logic_vector(13 downto 0);  -- rsp_xbar_mux_001:src_channel -> nios2_qsys_grms_data_master_translator_avalon_universal_master_0_agent:rp_channel
	signal rsp_xbar_mux_001_src_ready                                                                             : std_logic;                      -- nios2_qsys_grms_data_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux_001:src_ready
	signal cmd_xbar_mux_src_endofpacket                                                                           : std_logic;                      -- cmd_xbar_mux:src_endofpacket -> nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_src_valid                                                                                 : std_logic;                      -- cmd_xbar_mux:src_valid -> nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_src_startofpacket                                                                         : std_logic;                      -- cmd_xbar_mux:src_startofpacket -> nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_src_data                                                                                  : std_logic_vector(99 downto 0);  -- cmd_xbar_mux:src_data -> nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_src_channel                                                                               : std_logic_vector(13 downto 0);  -- cmd_xbar_mux:src_channel -> nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_src_ready                                                                                 : std_logic;                      -- nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	signal id_router_src_endofpacket                                                                              : std_logic;                      -- id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	signal id_router_src_valid                                                                                    : std_logic;                      -- id_router:src_valid -> rsp_xbar_demux:sink_valid
	signal id_router_src_startofpacket                                                                            : std_logic;                      -- id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	signal id_router_src_data                                                                                     : std_logic_vector(99 downto 0);  -- id_router:src_data -> rsp_xbar_demux:sink_data
	signal id_router_src_channel                                                                                  : std_logic_vector(13 downto 0);  -- id_router:src_channel -> rsp_xbar_demux:sink_channel
	signal id_router_src_ready                                                                                    : std_logic;                      -- rsp_xbar_demux:sink_ready -> id_router:src_ready
	signal cmd_xbar_mux_001_src_endofpacket                                                                       : std_logic;                      -- cmd_xbar_mux_001:src_endofpacket -> jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_001_src_valid                                                                             : std_logic;                      -- cmd_xbar_mux_001:src_valid -> jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_001_src_startofpacket                                                                     : std_logic;                      -- cmd_xbar_mux_001:src_startofpacket -> jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_001_src_data                                                                              : std_logic_vector(99 downto 0);  -- cmd_xbar_mux_001:src_data -> jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_001_src_channel                                                                           : std_logic_vector(13 downto 0);  -- cmd_xbar_mux_001:src_channel -> jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_001_src_ready                                                                             : std_logic;                      -- jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_001:src_ready
	signal id_router_001_src_endofpacket                                                                          : std_logic;                      -- id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	signal id_router_001_src_valid                                                                                : std_logic;                      -- id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	signal id_router_001_src_startofpacket                                                                        : std_logic;                      -- id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	signal id_router_001_src_data                                                                                 : std_logic_vector(99 downto 0);  -- id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	signal id_router_001_src_channel                                                                              : std_logic_vector(13 downto 0);  -- id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	signal id_router_001_src_ready                                                                                : std_logic;                      -- rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	signal cmd_xbar_mux_003_src_endofpacket                                                                       : std_logic;                      -- cmd_xbar_mux_003:src_endofpacket -> timer_grms_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_003_src_valid                                                                             : std_logic;                      -- cmd_xbar_mux_003:src_valid -> timer_grms_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_003_src_startofpacket                                                                     : std_logic;                      -- cmd_xbar_mux_003:src_startofpacket -> timer_grms_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_003_src_data                                                                              : std_logic_vector(99 downto 0);  -- cmd_xbar_mux_003:src_data -> timer_grms_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_003_src_channel                                                                           : std_logic_vector(13 downto 0);  -- cmd_xbar_mux_003:src_channel -> timer_grms_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_003_src_ready                                                                             : std_logic;                      -- timer_grms_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_003:src_ready
	signal id_router_003_src_endofpacket                                                                          : std_logic;                      -- id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	signal id_router_003_src_valid                                                                                : std_logic;                      -- id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	signal id_router_003_src_startofpacket                                                                        : std_logic;                      -- id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	signal id_router_003_src_data                                                                                 : std_logic_vector(99 downto 0);  -- id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	signal id_router_003_src_channel                                                                              : std_logic_vector(13 downto 0);  -- id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	signal id_router_003_src_ready                                                                                : std_logic;                      -- rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	signal cmd_xbar_mux_004_src_endofpacket                                                                       : std_logic;                      -- cmd_xbar_mux_004:src_endofpacket -> lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_004_src_valid                                                                             : std_logic;                      -- cmd_xbar_mux_004:src_valid -> lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_004_src_startofpacket                                                                     : std_logic;                      -- cmd_xbar_mux_004:src_startofpacket -> lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_004_src_data                                                                              : std_logic_vector(99 downto 0);  -- cmd_xbar_mux_004:src_data -> lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_004_src_channel                                                                           : std_logic_vector(13 downto 0);  -- cmd_xbar_mux_004:src_channel -> lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_004_src_ready                                                                             : std_logic;                      -- lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_004:src_ready
	signal id_router_004_src_endofpacket                                                                          : std_logic;                      -- id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	signal id_router_004_src_valid                                                                                : std_logic;                      -- id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	signal id_router_004_src_startofpacket                                                                        : std_logic;                      -- id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	signal id_router_004_src_data                                                                                 : std_logic_vector(99 downto 0);  -- id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	signal id_router_004_src_channel                                                                              : std_logic_vector(13 downto 0);  -- id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	signal id_router_004_src_ready                                                                                : std_logic;                      -- rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	signal cmd_xbar_mux_005_src_endofpacket                                                                       : std_logic;                      -- cmd_xbar_mux_005:src_endofpacket -> pa_grms_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_005_src_valid                                                                             : std_logic;                      -- cmd_xbar_mux_005:src_valid -> pa_grms_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_005_src_startofpacket                                                                     : std_logic;                      -- cmd_xbar_mux_005:src_startofpacket -> pa_grms_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_005_src_data                                                                              : std_logic_vector(99 downto 0);  -- cmd_xbar_mux_005:src_data -> pa_grms_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_005_src_channel                                                                           : std_logic_vector(13 downto 0);  -- cmd_xbar_mux_005:src_channel -> pa_grms_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_005_src_ready                                                                             : std_logic;                      -- pa_grms_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_005:src_ready
	signal id_router_005_src_endofpacket                                                                          : std_logic;                      -- id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	signal id_router_005_src_valid                                                                                : std_logic;                      -- id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	signal id_router_005_src_startofpacket                                                                        : std_logic;                      -- id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	signal id_router_005_src_data                                                                                 : std_logic_vector(99 downto 0);  -- id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	signal id_router_005_src_channel                                                                              : std_logic_vector(13 downto 0);  -- id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	signal id_router_005_src_ready                                                                                : std_logic;                      -- rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	signal cmd_xbar_mux_006_src_endofpacket                                                                       : std_logic;                      -- cmd_xbar_mux_006:src_endofpacket -> pb_grms_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_006_src_valid                                                                             : std_logic;                      -- cmd_xbar_mux_006:src_valid -> pb_grms_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_006_src_startofpacket                                                                     : std_logic;                      -- cmd_xbar_mux_006:src_startofpacket -> pb_grms_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_006_src_data                                                                              : std_logic_vector(99 downto 0);  -- cmd_xbar_mux_006:src_data -> pb_grms_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_006_src_channel                                                                           : std_logic_vector(13 downto 0);  -- cmd_xbar_mux_006:src_channel -> pb_grms_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_006_src_ready                                                                             : std_logic;                      -- pb_grms_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_006:src_ready
	signal id_router_006_src_endofpacket                                                                          : std_logic;                      -- id_router_006:src_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	signal id_router_006_src_valid                                                                                : std_logic;                      -- id_router_006:src_valid -> rsp_xbar_demux_006:sink_valid
	signal id_router_006_src_startofpacket                                                                        : std_logic;                      -- id_router_006:src_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	signal id_router_006_src_data                                                                                 : std_logic_vector(99 downto 0);  -- id_router_006:src_data -> rsp_xbar_demux_006:sink_data
	signal id_router_006_src_channel                                                                              : std_logic_vector(13 downto 0);  -- id_router_006:src_channel -> rsp_xbar_demux_006:sink_channel
	signal id_router_006_src_ready                                                                                : std_logic;                      -- rsp_xbar_demux_006:sink_ready -> id_router_006:src_ready
	signal cmd_xbar_mux_007_src_endofpacket                                                                       : std_logic;                      -- cmd_xbar_mux_007:src_endofpacket -> pc_grms_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_007_src_valid                                                                             : std_logic;                      -- cmd_xbar_mux_007:src_valid -> pc_grms_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_007_src_startofpacket                                                                     : std_logic;                      -- cmd_xbar_mux_007:src_startofpacket -> pc_grms_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_007_src_data                                                                              : std_logic_vector(99 downto 0);  -- cmd_xbar_mux_007:src_data -> pc_grms_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_007_src_channel                                                                           : std_logic_vector(13 downto 0);  -- cmd_xbar_mux_007:src_channel -> pc_grms_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_007_src_ready                                                                             : std_logic;                      -- pc_grms_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_007:src_ready
	signal id_router_007_src_endofpacket                                                                          : std_logic;                      -- id_router_007:src_endofpacket -> rsp_xbar_demux_007:sink_endofpacket
	signal id_router_007_src_valid                                                                                : std_logic;                      -- id_router_007:src_valid -> rsp_xbar_demux_007:sink_valid
	signal id_router_007_src_startofpacket                                                                        : std_logic;                      -- id_router_007:src_startofpacket -> rsp_xbar_demux_007:sink_startofpacket
	signal id_router_007_src_data                                                                                 : std_logic_vector(99 downto 0);  -- id_router_007:src_data -> rsp_xbar_demux_007:sink_data
	signal id_router_007_src_channel                                                                              : std_logic_vector(13 downto 0);  -- id_router_007:src_channel -> rsp_xbar_demux_007:sink_channel
	signal id_router_007_src_ready                                                                                : std_logic;                      -- rsp_xbar_demux_007:sink_ready -> id_router_007:src_ready
	signal cmd_xbar_mux_008_src_endofpacket                                                                       : std_logic;                      -- cmd_xbar_mux_008:src_endofpacket -> pd_grms_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_008_src_valid                                                                             : std_logic;                      -- cmd_xbar_mux_008:src_valid -> pd_grms_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_008_src_startofpacket                                                                     : std_logic;                      -- cmd_xbar_mux_008:src_startofpacket -> pd_grms_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_008_src_data                                                                              : std_logic_vector(99 downto 0);  -- cmd_xbar_mux_008:src_data -> pd_grms_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_008_src_channel                                                                           : std_logic_vector(13 downto 0);  -- cmd_xbar_mux_008:src_channel -> pd_grms_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_008_src_ready                                                                             : std_logic;                      -- pd_grms_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_008:src_ready
	signal id_router_008_src_endofpacket                                                                          : std_logic;                      -- id_router_008:src_endofpacket -> rsp_xbar_demux_008:sink_endofpacket
	signal id_router_008_src_valid                                                                                : std_logic;                      -- id_router_008:src_valid -> rsp_xbar_demux_008:sink_valid
	signal id_router_008_src_startofpacket                                                                        : std_logic;                      -- id_router_008:src_startofpacket -> rsp_xbar_demux_008:sink_startofpacket
	signal id_router_008_src_data                                                                                 : std_logic_vector(99 downto 0);  -- id_router_008:src_data -> rsp_xbar_demux_008:sink_data
	signal id_router_008_src_channel                                                                              : std_logic_vector(13 downto 0);  -- id_router_008:src_channel -> rsp_xbar_demux_008:sink_channel
	signal id_router_008_src_ready                                                                                : std_logic;                      -- rsp_xbar_demux_008:sink_ready -> id_router_008:src_ready
	signal cmd_xbar_mux_009_src_endofpacket                                                                       : std_logic;                      -- cmd_xbar_mux_009:src_endofpacket -> pe_grms_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_009_src_valid                                                                             : std_logic;                      -- cmd_xbar_mux_009:src_valid -> pe_grms_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_009_src_startofpacket                                                                     : std_logic;                      -- cmd_xbar_mux_009:src_startofpacket -> pe_grms_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_009_src_data                                                                              : std_logic_vector(99 downto 0);  -- cmd_xbar_mux_009:src_data -> pe_grms_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_009_src_channel                                                                           : std_logic_vector(13 downto 0);  -- cmd_xbar_mux_009:src_channel -> pe_grms_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_009_src_ready                                                                             : std_logic;                      -- pe_grms_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_009:src_ready
	signal id_router_009_src_endofpacket                                                                          : std_logic;                      -- id_router_009:src_endofpacket -> rsp_xbar_demux_009:sink_endofpacket
	signal id_router_009_src_valid                                                                                : std_logic;                      -- id_router_009:src_valid -> rsp_xbar_demux_009:sink_valid
	signal id_router_009_src_startofpacket                                                                        : std_logic;                      -- id_router_009:src_startofpacket -> rsp_xbar_demux_009:sink_startofpacket
	signal id_router_009_src_data                                                                                 : std_logic_vector(99 downto 0);  -- id_router_009:src_data -> rsp_xbar_demux_009:sink_data
	signal id_router_009_src_channel                                                                              : std_logic_vector(13 downto 0);  -- id_router_009:src_channel -> rsp_xbar_demux_009:sink_channel
	signal id_router_009_src_ready                                                                                : std_logic;                      -- rsp_xbar_demux_009:sink_ready -> id_router_009:src_ready
	signal cmd_xbar_mux_010_src_endofpacket                                                                       : std_logic;                      -- cmd_xbar_mux_010:src_endofpacket -> pf_grms_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_010_src_valid                                                                             : std_logic;                      -- cmd_xbar_mux_010:src_valid -> pf_grms_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_010_src_startofpacket                                                                     : std_logic;                      -- cmd_xbar_mux_010:src_startofpacket -> pf_grms_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_010_src_data                                                                              : std_logic_vector(99 downto 0);  -- cmd_xbar_mux_010:src_data -> pf_grms_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_010_src_channel                                                                           : std_logic_vector(13 downto 0);  -- cmd_xbar_mux_010:src_channel -> pf_grms_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_010_src_ready                                                                             : std_logic;                      -- pf_grms_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_010:src_ready
	signal id_router_010_src_endofpacket                                                                          : std_logic;                      -- id_router_010:src_endofpacket -> rsp_xbar_demux_010:sink_endofpacket
	signal id_router_010_src_valid                                                                                : std_logic;                      -- id_router_010:src_valid -> rsp_xbar_demux_010:sink_valid
	signal id_router_010_src_startofpacket                                                                        : std_logic;                      -- id_router_010:src_startofpacket -> rsp_xbar_demux_010:sink_startofpacket
	signal id_router_010_src_data                                                                                 : std_logic_vector(99 downto 0);  -- id_router_010:src_data -> rsp_xbar_demux_010:sink_data
	signal id_router_010_src_channel                                                                              : std_logic_vector(13 downto 0);  -- id_router_010:src_channel -> rsp_xbar_demux_010:sink_channel
	signal id_router_010_src_ready                                                                                : std_logic;                      -- rsp_xbar_demux_010:sink_ready -> id_router_010:src_ready
	signal cmd_xbar_mux_011_src_endofpacket                                                                       : std_logic;                      -- cmd_xbar_mux_011:src_endofpacket -> pg_grms_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_011_src_valid                                                                             : std_logic;                      -- cmd_xbar_mux_011:src_valid -> pg_grms_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_011_src_startofpacket                                                                     : std_logic;                      -- cmd_xbar_mux_011:src_startofpacket -> pg_grms_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_011_src_data                                                                              : std_logic_vector(99 downto 0);  -- cmd_xbar_mux_011:src_data -> pg_grms_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_011_src_channel                                                                           : std_logic_vector(13 downto 0);  -- cmd_xbar_mux_011:src_channel -> pg_grms_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_011_src_ready                                                                             : std_logic;                      -- pg_grms_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_011:src_ready
	signal id_router_011_src_endofpacket                                                                          : std_logic;                      -- id_router_011:src_endofpacket -> rsp_xbar_demux_011:sink_endofpacket
	signal id_router_011_src_valid                                                                                : std_logic;                      -- id_router_011:src_valid -> rsp_xbar_demux_011:sink_valid
	signal id_router_011_src_startofpacket                                                                        : std_logic;                      -- id_router_011:src_startofpacket -> rsp_xbar_demux_011:sink_startofpacket
	signal id_router_011_src_data                                                                                 : std_logic_vector(99 downto 0);  -- id_router_011:src_data -> rsp_xbar_demux_011:sink_data
	signal id_router_011_src_channel                                                                              : std_logic_vector(13 downto 0);  -- id_router_011:src_channel -> rsp_xbar_demux_011:sink_channel
	signal id_router_011_src_ready                                                                                : std_logic;                      -- rsp_xbar_demux_011:sink_ready -> id_router_011:src_ready
	signal cmd_xbar_mux_012_src_endofpacket                                                                       : std_logic;                      -- cmd_xbar_mux_012:src_endofpacket -> ph_grms_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_012_src_valid                                                                             : std_logic;                      -- cmd_xbar_mux_012:src_valid -> ph_grms_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_012_src_startofpacket                                                                     : std_logic;                      -- cmd_xbar_mux_012:src_startofpacket -> ph_grms_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_012_src_data                                                                              : std_logic_vector(99 downto 0);  -- cmd_xbar_mux_012:src_data -> ph_grms_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_012_src_channel                                                                           : std_logic_vector(13 downto 0);  -- cmd_xbar_mux_012:src_channel -> ph_grms_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_012_src_ready                                                                             : std_logic;                      -- ph_grms_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_012:src_ready
	signal id_router_012_src_endofpacket                                                                          : std_logic;                      -- id_router_012:src_endofpacket -> rsp_xbar_demux_012:sink_endofpacket
	signal id_router_012_src_valid                                                                                : std_logic;                      -- id_router_012:src_valid -> rsp_xbar_demux_012:sink_valid
	signal id_router_012_src_startofpacket                                                                        : std_logic;                      -- id_router_012:src_startofpacket -> rsp_xbar_demux_012:sink_startofpacket
	signal id_router_012_src_data                                                                                 : std_logic_vector(99 downto 0);  -- id_router_012:src_data -> rsp_xbar_demux_012:sink_data
	signal id_router_012_src_channel                                                                              : std_logic_vector(13 downto 0);  -- id_router_012:src_channel -> rsp_xbar_demux_012:sink_channel
	signal id_router_012_src_ready                                                                                : std_logic;                      -- rsp_xbar_demux_012:sink_ready -> id_router_012:src_ready
	signal cmd_xbar_mux_013_src_endofpacket                                                                       : std_logic;                      -- cmd_xbar_mux_013:src_endofpacket -> pi_grms_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_013_src_valid                                                                             : std_logic;                      -- cmd_xbar_mux_013:src_valid -> pi_grms_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_013_src_startofpacket                                                                     : std_logic;                      -- cmd_xbar_mux_013:src_startofpacket -> pi_grms_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_013_src_data                                                                              : std_logic_vector(99 downto 0);  -- cmd_xbar_mux_013:src_data -> pi_grms_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_013_src_channel                                                                           : std_logic_vector(13 downto 0);  -- cmd_xbar_mux_013:src_channel -> pi_grms_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_013_src_ready                                                                             : std_logic;                      -- pi_grms_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_013:src_ready
	signal id_router_013_src_endofpacket                                                                          : std_logic;                      -- id_router_013:src_endofpacket -> rsp_xbar_demux_013:sink_endofpacket
	signal id_router_013_src_valid                                                                                : std_logic;                      -- id_router_013:src_valid -> rsp_xbar_demux_013:sink_valid
	signal id_router_013_src_startofpacket                                                                        : std_logic;                      -- id_router_013:src_startofpacket -> rsp_xbar_demux_013:sink_startofpacket
	signal id_router_013_src_data                                                                                 : std_logic_vector(99 downto 0);  -- id_router_013:src_data -> rsp_xbar_demux_013:sink_data
	signal id_router_013_src_channel                                                                              : std_logic_vector(13 downto 0);  -- id_router_013:src_channel -> rsp_xbar_demux_013:sink_channel
	signal id_router_013_src_ready                                                                                : std_logic;                      -- rsp_xbar_demux_013:sink_ready -> id_router_013:src_ready
	signal cmd_xbar_mux_002_src_endofpacket                                                                       : std_logic;                      -- cmd_xbar_mux_002:src_endofpacket -> width_adapter:in_endofpacket
	signal cmd_xbar_mux_002_src_valid                                                                             : std_logic;                      -- cmd_xbar_mux_002:src_valid -> width_adapter:in_valid
	signal cmd_xbar_mux_002_src_startofpacket                                                                     : std_logic;                      -- cmd_xbar_mux_002:src_startofpacket -> width_adapter:in_startofpacket
	signal cmd_xbar_mux_002_src_data                                                                              : std_logic_vector(99 downto 0);  -- cmd_xbar_mux_002:src_data -> width_adapter:in_data
	signal cmd_xbar_mux_002_src_channel                                                                           : std_logic_vector(13 downto 0);  -- cmd_xbar_mux_002:src_channel -> width_adapter:in_channel
	signal cmd_xbar_mux_002_src_ready                                                                             : std_logic;                      -- width_adapter:in_ready -> cmd_xbar_mux_002:src_ready
	signal width_adapter_src_endofpacket                                                                          : std_logic;                      -- width_adapter:out_endofpacket -> burst_adapter:sink0_endofpacket
	signal width_adapter_src_valid                                                                                : std_logic;                      -- width_adapter:out_valid -> burst_adapter:sink0_valid
	signal width_adapter_src_startofpacket                                                                        : std_logic;                      -- width_adapter:out_startofpacket -> burst_adapter:sink0_startofpacket
	signal width_adapter_src_data                                                                                 : std_logic_vector(81 downto 0);  -- width_adapter:out_data -> burst_adapter:sink0_data
	signal width_adapter_src_ready                                                                                : std_logic;                      -- burst_adapter:sink0_ready -> width_adapter:out_ready
	signal width_adapter_src_channel                                                                              : std_logic_vector(13 downto 0);  -- width_adapter:out_channel -> burst_adapter:sink0_channel
	signal id_router_002_src_endofpacket                                                                          : std_logic;                      -- id_router_002:src_endofpacket -> width_adapter_001:in_endofpacket
	signal id_router_002_src_valid                                                                                : std_logic;                      -- id_router_002:src_valid -> width_adapter_001:in_valid
	signal id_router_002_src_startofpacket                                                                        : std_logic;                      -- id_router_002:src_startofpacket -> width_adapter_001:in_startofpacket
	signal id_router_002_src_data                                                                                 : std_logic_vector(81 downto 0);  -- id_router_002:src_data -> width_adapter_001:in_data
	signal id_router_002_src_channel                                                                              : std_logic_vector(13 downto 0);  -- id_router_002:src_channel -> width_adapter_001:in_channel
	signal id_router_002_src_ready                                                                                : std_logic;                      -- width_adapter_001:in_ready -> id_router_002:src_ready
	signal width_adapter_001_src_endofpacket                                                                      : std_logic;                      -- width_adapter_001:out_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	signal width_adapter_001_src_valid                                                                            : std_logic;                      -- width_adapter_001:out_valid -> rsp_xbar_demux_002:sink_valid
	signal width_adapter_001_src_startofpacket                                                                    : std_logic;                      -- width_adapter_001:out_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	signal width_adapter_001_src_data                                                                             : std_logic_vector(99 downto 0);  -- width_adapter_001:out_data -> rsp_xbar_demux_002:sink_data
	signal width_adapter_001_src_ready                                                                            : std_logic;                      -- rsp_xbar_demux_002:sink_ready -> width_adapter_001:out_ready
	signal width_adapter_001_src_channel                                                                          : std_logic_vector(13 downto 0);  -- width_adapter_001:out_channel -> rsp_xbar_demux_002:sink_channel
	signal irq_mapper_receiver0_irq                                                                               : std_logic;                      -- jtag_uart_grms:av_irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                                                               : std_logic;                      -- timer_grms:irq -> irq_mapper:receiver1_irq
	signal nios2_qsys_grms_d_irq_irq                                                                              : std_logic_vector(31 downto 0);  -- irq_mapper:sender_irq -> nios2_qsys_grms:d_irq
	signal reset_reset_n_ports_inv                                                                                : std_logic;                      -- reset_reset_n:inv -> rst_controller:reset_in0
	signal jtag_uart_grms_avalon_jtag_slave_translator_avalon_anti_slave_0_write_ports_inv                        : std_logic;                      -- jtag_uart_grms_avalon_jtag_slave_translator_avalon_anti_slave_0_write:inv -> jtag_uart_grms:av_write_n
	signal jtag_uart_grms_avalon_jtag_slave_translator_avalon_anti_slave_0_read_ports_inv                         : std_logic;                      -- jtag_uart_grms_avalon_jtag_slave_translator_avalon_anti_slave_0_read:inv -> jtag_uart_grms:av_read_n
	signal new_sdram_controller_grms_s1_translator_avalon_anti_slave_0_write_ports_inv                            : std_logic;                      -- new_sdram_controller_grms_s1_translator_avalon_anti_slave_0_write:inv -> new_sdram_controller_grms:az_wr_n
	signal new_sdram_controller_grms_s1_translator_avalon_anti_slave_0_read_ports_inv                             : std_logic;                      -- new_sdram_controller_grms_s1_translator_avalon_anti_slave_0_read:inv -> new_sdram_controller_grms:az_rd_n
	signal new_sdram_controller_grms_s1_translator_avalon_anti_slave_0_byteenable_ports_inv                       : std_logic_vector(1 downto 0);   -- new_sdram_controller_grms_s1_translator_avalon_anti_slave_0_byteenable:inv -> new_sdram_controller_grms:az_be_n
	signal timer_grms_s1_translator_avalon_anti_slave_0_write_ports_inv                                           : std_logic;                      -- timer_grms_s1_translator_avalon_anti_slave_0_write:inv -> timer_grms:write_n
	signal pc_grms_s1_translator_avalon_anti_slave_0_write_ports_inv                                              : std_logic;                      -- pc_grms_s1_translator_avalon_anti_slave_0_write:inv -> pc_grms:write_n
	signal pd_grms_s1_translator_avalon_anti_slave_0_write_ports_inv                                              : std_logic;                      -- pd_grms_s1_translator_avalon_anti_slave_0_write:inv -> pd_grms:write_n
	signal pe_grms_s1_translator_avalon_anti_slave_0_write_ports_inv                                              : std_logic;                      -- pe_grms_s1_translator_avalon_anti_slave_0_write:inv -> pe_grms:write_n
	signal pf_grms_s1_translator_avalon_anti_slave_0_write_ports_inv                                              : std_logic;                      -- pf_grms_s1_translator_avalon_anti_slave_0_write:inv -> pf_grms:write_n
	signal pg_grms_s1_translator_avalon_anti_slave_0_write_ports_inv                                              : std_logic;                      -- pg_grms_s1_translator_avalon_anti_slave_0_write:inv -> pg_grms:write_n
	signal ph_grms_s1_translator_avalon_anti_slave_0_write_ports_inv                                              : std_logic;                      -- ph_grms_s1_translator_avalon_anti_slave_0_write:inv -> ph_grms:write_n
	signal pi_grms_s1_translator_avalon_anti_slave_0_write_ports_inv                                              : std_logic;                      -- pi_grms_s1_translator_avalon_anti_slave_0_write:inv -> pi_grms:write_n
	signal rst_controller_reset_out_reset_ports_inv                                                               : std_logic;                      -- rst_controller_reset_out_reset:inv -> [jtag_uart_grms:rst_n, lcd_16207_grms:reset_n, new_sdram_controller_grms:reset_n, nios2_qsys_grms:reset_n, pa_grms:reset_n, pb_grms:reset_n, pc_grms:reset_n, pd_grms:reset_n, pe_grms:reset_n, pf_grms:reset_n, pg_grms:reset_n, ph_grms:reset_n, pi_grms:reset_n, timer_grms:reset_n]

begin

	nios2_qsys_grms : component p2_grms_qsys_nios2_qsys_grms
		port map (
			clk                                   => clk_clk,                                                                      --                       clk.clk
			reset_n                               => rst_controller_reset_out_reset_ports_inv,                                     --                   reset_n.reset_n
			d_address                             => nios2_qsys_grms_data_master_address,                                          --               data_master.address
			d_byteenable                          => nios2_qsys_grms_data_master_byteenable,                                       --                          .byteenable
			d_read                                => nios2_qsys_grms_data_master_read,                                             --                          .read
			d_readdata                            => nios2_qsys_grms_data_master_readdata,                                         --                          .readdata
			d_waitrequest                         => nios2_qsys_grms_data_master_waitrequest,                                      --                          .waitrequest
			d_write                               => nios2_qsys_grms_data_master_write,                                            --                          .write
			d_writedata                           => nios2_qsys_grms_data_master_writedata,                                        --                          .writedata
			jtag_debug_module_debugaccess_to_roms => nios2_qsys_grms_data_master_debugaccess,                                      --                          .debugaccess
			i_address                             => nios2_qsys_grms_instruction_master_address,                                   --        instruction_master.address
			i_read                                => nios2_qsys_grms_instruction_master_read,                                      --                          .read
			i_readdata                            => nios2_qsys_grms_instruction_master_readdata,                                  --                          .readdata
			i_waitrequest                         => nios2_qsys_grms_instruction_master_waitrequest,                               --                          .waitrequest
			d_irq                                 => nios2_qsys_grms_d_irq_irq,                                                    --                     d_irq.irq
			jtag_debug_module_resetrequest        => open,                                                                         --   jtag_debug_module_reset.reset
			jtag_debug_module_address             => nios2_qsys_grms_jtag_debug_module_translator_avalon_anti_slave_0_address,     --         jtag_debug_module.address
			jtag_debug_module_byteenable          => nios2_qsys_grms_jtag_debug_module_translator_avalon_anti_slave_0_byteenable,  --                          .byteenable
			jtag_debug_module_debugaccess         => nios2_qsys_grms_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess, --                          .debugaccess
			jtag_debug_module_read                => nios2_qsys_grms_jtag_debug_module_translator_avalon_anti_slave_0_read,        --                          .read
			jtag_debug_module_readdata            => nios2_qsys_grms_jtag_debug_module_translator_avalon_anti_slave_0_readdata,    --                          .readdata
			jtag_debug_module_waitrequest         => nios2_qsys_grms_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest, --                          .waitrequest
			jtag_debug_module_write               => nios2_qsys_grms_jtag_debug_module_translator_avalon_anti_slave_0_write,       --                          .write
			jtag_debug_module_writedata           => nios2_qsys_grms_jtag_debug_module_translator_avalon_anti_slave_0_writedata,   --                          .writedata
			no_ci_readra                          => open                                                                          -- custom_instruction_master.readra
		);

	jtag_uart_grms : component p2_grms_qsys_jtag_uart_grms
		port map (
			clk            => clk_clk,                                                                         --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                                        --             reset.reset_n
			av_chipselect  => jtag_uart_grms_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => jtag_uart_grms_avalon_jtag_slave_translator_avalon_anti_slave_0_address(0),      --                  .address
			av_read_n      => jtag_uart_grms_avalon_jtag_slave_translator_avalon_anti_slave_0_read_ports_inv,  --                  .read_n
			av_readdata    => jtag_uart_grms_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata,        --                  .readdata
			av_write_n     => jtag_uart_grms_avalon_jtag_slave_translator_avalon_anti_slave_0_write_ports_inv, --                  .write_n
			av_writedata   => jtag_uart_grms_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata,       --                  .writedata
			av_waitrequest => jtag_uart_grms_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver0_irq                                                         --               irq.irq
		);

	new_sdram_controller_grms : component p2_grms_qsys_new_sdram_controller_grms
		port map (
			clk            => clk_clk,                                                                          --   clk.clk
			reset_n        => rst_controller_reset_out_reset_ports_inv,                                         -- reset.reset_n
			az_addr        => new_sdram_controller_grms_s1_translator_avalon_anti_slave_0_address,              --    s1.address
			az_be_n        => new_sdram_controller_grms_s1_translator_avalon_anti_slave_0_byteenable_ports_inv, --      .byteenable_n
			az_cs          => new_sdram_controller_grms_s1_translator_avalon_anti_slave_0_chipselect,           --      .chipselect
			az_data        => new_sdram_controller_grms_s1_translator_avalon_anti_slave_0_writedata,            --      .writedata
			az_rd_n        => new_sdram_controller_grms_s1_translator_avalon_anti_slave_0_read_ports_inv,       --      .read_n
			az_wr_n        => new_sdram_controller_grms_s1_translator_avalon_anti_slave_0_write_ports_inv,      --      .write_n
			za_data        => new_sdram_controller_grms_s1_translator_avalon_anti_slave_0_readdata,             --      .readdata
			za_valid       => new_sdram_controller_grms_s1_translator_avalon_anti_slave_0_readdatavalid,        --      .readdatavalid
			za_waitrequest => new_sdram_controller_grms_s1_translator_avalon_anti_slave_0_waitrequest,          --      .waitrequest
			zs_addr        => new_sdram_controller_grms_wire_addr,                                              --  wire.export
			zs_ba          => new_sdram_controller_grms_wire_ba,                                                --      .export
			zs_cas_n       => new_sdram_controller_grms_wire_cas_n,                                             --      .export
			zs_cke         => new_sdram_controller_grms_wire_cke,                                               --      .export
			zs_cs_n        => new_sdram_controller_grms_wire_cs_n,                                              --      .export
			zs_dq          => new_sdram_controller_grms_wire_dq,                                                --      .export
			zs_dqm         => new_sdram_controller_grms_wire_dqm,                                               --      .export
			zs_ras_n       => new_sdram_controller_grms_wire_ras_n,                                             --      .export
			zs_we_n        => new_sdram_controller_grms_wire_we_n                                               --      .export
		);

	timer_grms : component p2_grms_qsys_timer_grms
		port map (
			clk        => clk_clk,                                                      --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                     -- reset.reset_n
			address    => timer_grms_s1_translator_avalon_anti_slave_0_address,         --    s1.address
			writedata  => timer_grms_s1_translator_avalon_anti_slave_0_writedata,       --      .writedata
			readdata   => timer_grms_s1_translator_avalon_anti_slave_0_readdata,        --      .readdata
			chipselect => timer_grms_s1_translator_avalon_anti_slave_0_chipselect,      --      .chipselect
			write_n    => timer_grms_s1_translator_avalon_anti_slave_0_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver1_irq                                      --   irq.irq
		);

	lcd_16207_grms : component p2_grms_qsys_lcd_16207_grms
		port map (
			reset_n       => rst_controller_reset_out_reset_ports_inv,                                  --         reset.reset_n
			clk           => clk_clk,                                                                   --           clk.clk
			begintransfer => lcd_16207_grms_control_slave_translator_avalon_anti_slave_0_begintransfer, -- control_slave.begintransfer
			read          => lcd_16207_grms_control_slave_translator_avalon_anti_slave_0_read,          --              .read
			write         => lcd_16207_grms_control_slave_translator_avalon_anti_slave_0_write,         --              .write
			readdata      => lcd_16207_grms_control_slave_translator_avalon_anti_slave_0_readdata,      --              .readdata
			writedata     => lcd_16207_grms_control_slave_translator_avalon_anti_slave_0_writedata,     --              .writedata
			address       => lcd_16207_grms_control_slave_translator_avalon_anti_slave_0_address,       --              .address
			LCD_RS        => lcd_16207_grms_external_RS,                                                --      external.export
			LCD_RW        => lcd_16207_grms_external_RW,                                                --              .export
			LCD_data      => lcd_16207_grms_external_data,                                              --              .export
			LCD_E         => lcd_16207_grms_external_E                                                  --              .export
		);

	pa_grms : component p2_grms_qsys_pa_grms
		port map (
			clk      => clk_clk,                                            --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,           --               reset.reset_n
			address  => pa_grms_s1_translator_avalon_anti_slave_0_address,  --                  s1.address
			readdata => pa_grms_s1_translator_avalon_anti_slave_0_readdata, --                    .readdata
			in_port  => pa_grms_external_connection_export                  -- external_connection.export
		);

	pb_grms : component p2_grms_qsys_pb_grms
		port map (
			clk      => clk_clk,                                            --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,           --               reset.reset_n
			address  => pb_grms_s1_translator_avalon_anti_slave_0_address,  --                  s1.address
			readdata => pb_grms_s1_translator_avalon_anti_slave_0_readdata, --                    .readdata
			in_port  => pb_grms_external_connection_export                  -- external_connection.export
		);

	pc_grms : component p2_grms_qsys_pc_grms
		port map (
			clk        => clk_clk,                                                   --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                  --               reset.reset_n
			address    => pc_grms_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => pc_grms_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => pc_grms_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => pc_grms_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => pc_grms_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			out_port   => pc_grms_external_connection_export                         -- external_connection.export
		);

	pd_grms : component p2_grms_qsys_pd_grms
		port map (
			clk        => clk_clk,                                                   --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                  --               reset.reset_n
			address    => pd_grms_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => pd_grms_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => pd_grms_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => pd_grms_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => pd_grms_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			out_port   => pd_grms_external_connection_export                         -- external_connection.export
		);

	pe_grms : component p2_grms_qsys_pd_grms
		port map (
			clk        => clk_clk,                                                   --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                  --               reset.reset_n
			address    => pe_grms_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => pe_grms_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => pe_grms_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => pe_grms_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => pe_grms_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			out_port   => pe_grms_external_connection_export                         -- external_connection.export
		);

	pf_grms : component p2_grms_qsys_pf_grms
		port map (
			clk        => clk_clk,                                                   --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                  --               reset.reset_n
			address    => pf_grms_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => pf_grms_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => pf_grms_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => pf_grms_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => pf_grms_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			out_port   => pf_grms_external_connection_export                         -- external_connection.export
		);

	pg_grms : component p2_grms_qsys_pf_grms
		port map (
			clk        => clk_clk,                                                   --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                  --               reset.reset_n
			address    => pg_grms_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => pg_grms_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => pg_grms_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => pg_grms_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => pg_grms_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			out_port   => pg_grms_external_connection_export                         -- external_connection.export
		);

	ph_grms : component p2_grms_qsys_ph_grms
		port map (
			clk        => clk_clk,                                                   --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                  --               reset.reset_n
			address    => ph_grms_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => ph_grms_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => ph_grms_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => ph_grms_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => ph_grms_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			out_port   => ph_grms_external_connection_export                         -- external_connection.export
		);

	pi_grms : component p2_grms_qsys_ph_grms
		port map (
			clk        => clk_clk,                                                   --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                  --               reset.reset_n
			address    => pi_grms_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => pi_grms_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => pi_grms_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => pi_grms_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => pi_grms_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			out_port   => pi_grms_external_connection_export                         -- external_connection.export
		);

	nios2_qsys_grms_instruction_master_translator : component p2_grms_qsys_nios2_qsys_grms_instruction_master_translator
		generic map (
			AV_ADDRESS_W                => 25,
			AV_DATA_W                   => 32,
			AV_BURSTCOUNT_W             => 1,
			AV_BYTEENABLE_W             => 4,
			UAV_ADDRESS_W               => 25,
			UAV_BURSTCOUNT_W            => 3,
			USE_READ                    => 1,
			USE_WRITE                   => 0,
			USE_BEGINBURSTTRANSFER      => 0,
			USE_BEGINTRANSFER           => 0,
			USE_CHIPSELECT              => 0,
			USE_BURSTCOUNT              => 0,
			USE_READDATAVALID           => 0,
			USE_WAITREQUEST             => 1,
			USE_READRESPONSE            => 0,
			USE_WRITERESPONSE           => 0,
			AV_SYMBOLS_PER_WORD         => 4,
			AV_ADDRESS_SYMBOLS          => 1,
			AV_BURSTCOUNT_SYMBOLS       => 0,
			AV_CONSTANT_BURST_BEHAVIOR  => 0,
			UAV_CONSTANT_BURST_BEHAVIOR => 0,
			AV_LINEWRAPBURSTS           => 1,
			AV_REGISTERINCOMINGSIGNALS  => 0
		)
		port map (
			clk                      => clk_clk,                                                                               --                       clk.clk
			reset                    => rst_controller_reset_out_reset,                                                        --                     reset.reset
			uav_address              => nios2_qsys_grms_instruction_master_translator_avalon_universal_master_0_address,       -- avalon_universal_master_0.address
			uav_burstcount           => nios2_qsys_grms_instruction_master_translator_avalon_universal_master_0_burstcount,    --                          .burstcount
			uav_read                 => nios2_qsys_grms_instruction_master_translator_avalon_universal_master_0_read,          --                          .read
			uav_write                => nios2_qsys_grms_instruction_master_translator_avalon_universal_master_0_write,         --                          .write
			uav_waitrequest          => nios2_qsys_grms_instruction_master_translator_avalon_universal_master_0_waitrequest,   --                          .waitrequest
			uav_readdatavalid        => nios2_qsys_grms_instruction_master_translator_avalon_universal_master_0_readdatavalid, --                          .readdatavalid
			uav_byteenable           => nios2_qsys_grms_instruction_master_translator_avalon_universal_master_0_byteenable,    --                          .byteenable
			uav_readdata             => nios2_qsys_grms_instruction_master_translator_avalon_universal_master_0_readdata,      --                          .readdata
			uav_writedata            => nios2_qsys_grms_instruction_master_translator_avalon_universal_master_0_writedata,     --                          .writedata
			uav_lock                 => nios2_qsys_grms_instruction_master_translator_avalon_universal_master_0_lock,          --                          .lock
			uav_debugaccess          => nios2_qsys_grms_instruction_master_translator_avalon_universal_master_0_debugaccess,   --                          .debugaccess
			av_address               => nios2_qsys_grms_instruction_master_address,                                            --      avalon_anti_master_0.address
			av_waitrequest           => nios2_qsys_grms_instruction_master_waitrequest,                                        --                          .waitrequest
			av_read                  => nios2_qsys_grms_instruction_master_read,                                               --                          .read
			av_readdata              => nios2_qsys_grms_instruction_master_readdata,                                           --                          .readdata
			av_burstcount            => "1",                                                                                   --               (terminated)
			av_byteenable            => "1111",                                                                                --               (terminated)
			av_beginbursttransfer    => '0',                                                                                   --               (terminated)
			av_begintransfer         => '0',                                                                                   --               (terminated)
			av_chipselect            => '0',                                                                                   --               (terminated)
			av_readdatavalid         => open,                                                                                  --               (terminated)
			av_write                 => '0',                                                                                   --               (terminated)
			av_writedata             => "00000000000000000000000000000000",                                                    --               (terminated)
			av_lock                  => '0',                                                                                   --               (terminated)
			av_debugaccess           => '0',                                                                                   --               (terminated)
			uav_clken                => open,                                                                                  --               (terminated)
			av_clken                 => '1',                                                                                   --               (terminated)
			uav_response             => "00",                                                                                  --               (terminated)
			av_response              => open,                                                                                  --               (terminated)
			uav_writeresponserequest => open,                                                                                  --               (terminated)
			uav_writeresponsevalid   => '0',                                                                                   --               (terminated)
			av_writeresponserequest  => '0',                                                                                   --               (terminated)
			av_writeresponsevalid    => open                                                                                   --               (terminated)
		);

	nios2_qsys_grms_data_master_translator : component p2_grms_qsys_nios2_qsys_grms_data_master_translator
		generic map (
			AV_ADDRESS_W                => 25,
			AV_DATA_W                   => 32,
			AV_BURSTCOUNT_W             => 1,
			AV_BYTEENABLE_W             => 4,
			UAV_ADDRESS_W               => 25,
			UAV_BURSTCOUNT_W            => 3,
			USE_READ                    => 1,
			USE_WRITE                   => 1,
			USE_BEGINBURSTTRANSFER      => 0,
			USE_BEGINTRANSFER           => 0,
			USE_CHIPSELECT              => 0,
			USE_BURSTCOUNT              => 0,
			USE_READDATAVALID           => 0,
			USE_WAITREQUEST             => 1,
			USE_READRESPONSE            => 0,
			USE_WRITERESPONSE           => 0,
			AV_SYMBOLS_PER_WORD         => 4,
			AV_ADDRESS_SYMBOLS          => 1,
			AV_BURSTCOUNT_SYMBOLS       => 0,
			AV_CONSTANT_BURST_BEHAVIOR  => 0,
			UAV_CONSTANT_BURST_BEHAVIOR => 0,
			AV_LINEWRAPBURSTS           => 0,
			AV_REGISTERINCOMINGSIGNALS  => 1
		)
		port map (
			clk                      => clk_clk,                                                                        --                       clk.clk
			reset                    => rst_controller_reset_out_reset,                                                 --                     reset.reset
			uav_address              => nios2_qsys_grms_data_master_translator_avalon_universal_master_0_address,       -- avalon_universal_master_0.address
			uav_burstcount           => nios2_qsys_grms_data_master_translator_avalon_universal_master_0_burstcount,    --                          .burstcount
			uav_read                 => nios2_qsys_grms_data_master_translator_avalon_universal_master_0_read,          --                          .read
			uav_write                => nios2_qsys_grms_data_master_translator_avalon_universal_master_0_write,         --                          .write
			uav_waitrequest          => nios2_qsys_grms_data_master_translator_avalon_universal_master_0_waitrequest,   --                          .waitrequest
			uav_readdatavalid        => nios2_qsys_grms_data_master_translator_avalon_universal_master_0_readdatavalid, --                          .readdatavalid
			uav_byteenable           => nios2_qsys_grms_data_master_translator_avalon_universal_master_0_byteenable,    --                          .byteenable
			uav_readdata             => nios2_qsys_grms_data_master_translator_avalon_universal_master_0_readdata,      --                          .readdata
			uav_writedata            => nios2_qsys_grms_data_master_translator_avalon_universal_master_0_writedata,     --                          .writedata
			uav_lock                 => nios2_qsys_grms_data_master_translator_avalon_universal_master_0_lock,          --                          .lock
			uav_debugaccess          => nios2_qsys_grms_data_master_translator_avalon_universal_master_0_debugaccess,   --                          .debugaccess
			av_address               => nios2_qsys_grms_data_master_address,                                            --      avalon_anti_master_0.address
			av_waitrequest           => nios2_qsys_grms_data_master_waitrequest,                                        --                          .waitrequest
			av_byteenable            => nios2_qsys_grms_data_master_byteenable,                                         --                          .byteenable
			av_read                  => nios2_qsys_grms_data_master_read,                                               --                          .read
			av_readdata              => nios2_qsys_grms_data_master_readdata,                                           --                          .readdata
			av_write                 => nios2_qsys_grms_data_master_write,                                              --                          .write
			av_writedata             => nios2_qsys_grms_data_master_writedata,                                          --                          .writedata
			av_debugaccess           => nios2_qsys_grms_data_master_debugaccess,                                        --                          .debugaccess
			av_burstcount            => "1",                                                                            --               (terminated)
			av_beginbursttransfer    => '0',                                                                            --               (terminated)
			av_begintransfer         => '0',                                                                            --               (terminated)
			av_chipselect            => '0',                                                                            --               (terminated)
			av_readdatavalid         => open,                                                                           --               (terminated)
			av_lock                  => '0',                                                                            --               (terminated)
			uav_clken                => open,                                                                           --               (terminated)
			av_clken                 => '1',                                                                            --               (terminated)
			uav_response             => "00",                                                                           --               (terminated)
			av_response              => open,                                                                           --               (terminated)
			uav_writeresponserequest => open,                                                                           --               (terminated)
			uav_writeresponsevalid   => '0',                                                                            --               (terminated)
			av_writeresponserequest  => '0',                                                                            --               (terminated)
			av_writeresponsevalid    => open                                                                            --               (terminated)
		);

	nios2_qsys_grms_jtag_debug_module_translator : component p2_grms_qsys_nios2_qsys_grms_jtag_debug_module_translator
		generic map (
			AV_ADDRESS_W                   => 9,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 1,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                                                      --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                               --                    reset.reset
			uav_address              => nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => nios2_qsys_grms_jtag_debug_module_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => nios2_qsys_grms_jtag_debug_module_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => nios2_qsys_grms_jtag_debug_module_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => nios2_qsys_grms_jtag_debug_module_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => nios2_qsys_grms_jtag_debug_module_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_byteenable            => nios2_qsys_grms_jtag_debug_module_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_waitrequest           => nios2_qsys_grms_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest,                 --                         .waitrequest
			av_debugaccess           => nios2_qsys_grms_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess,                 --                         .debugaccess
			av_begintransfer         => open,                                                                                         --              (terminated)
			av_beginbursttransfer    => open,                                                                                         --              (terminated)
			av_burstcount            => open,                                                                                         --              (terminated)
			av_readdatavalid         => '0',                                                                                          --              (terminated)
			av_writebyteenable       => open,                                                                                         --              (terminated)
			av_lock                  => open,                                                                                         --              (terminated)
			av_chipselect            => open,                                                                                         --              (terminated)
			av_clken                 => open,                                                                                         --              (terminated)
			uav_clken                => '0',                                                                                          --              (terminated)
			av_outputenable          => open,                                                                                         --              (terminated)
			uav_response             => open,                                                                                         --              (terminated)
			av_response              => "00",                                                                                         --              (terminated)
			uav_writeresponserequest => '0',                                                                                          --              (terminated)
			uav_writeresponsevalid   => open,                                                                                         --              (terminated)
			av_writeresponserequest  => open,                                                                                         --              (terminated)
			av_writeresponsevalid    => '0'                                                                                           --              (terminated)
		);

	jtag_uart_grms_avalon_jtag_slave_translator : component p2_grms_qsys_jtag_uart_grms_avalon_jtag_slave_translator
		generic map (
			AV_ADDRESS_W                   => 1,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 1,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                                                     --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                              --                    reset.reset
			uav_address              => jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => jtag_uart_grms_avalon_jtag_slave_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => jtag_uart_grms_avalon_jtag_slave_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => jtag_uart_grms_avalon_jtag_slave_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => jtag_uart_grms_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => jtag_uart_grms_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_waitrequest           => jtag_uart_grms_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest,                 --                         .waitrequest
			av_chipselect            => jtag_uart_grms_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_begintransfer         => open,                                                                                        --              (terminated)
			av_beginbursttransfer    => open,                                                                                        --              (terminated)
			av_burstcount            => open,                                                                                        --              (terminated)
			av_byteenable            => open,                                                                                        --              (terminated)
			av_readdatavalid         => '0',                                                                                         --              (terminated)
			av_writebyteenable       => open,                                                                                        --              (terminated)
			av_lock                  => open,                                                                                        --              (terminated)
			av_clken                 => open,                                                                                        --              (terminated)
			uav_clken                => '0',                                                                                         --              (terminated)
			av_debugaccess           => open,                                                                                        --              (terminated)
			av_outputenable          => open,                                                                                        --              (terminated)
			uav_response             => open,                                                                                        --              (terminated)
			av_response              => "00",                                                                                        --              (terminated)
			uav_writeresponserequest => '0',                                                                                         --              (terminated)
			uav_writeresponsevalid   => open,                                                                                        --              (terminated)
			av_writeresponserequest  => open,                                                                                        --              (terminated)
			av_writeresponsevalid    => '0'                                                                                          --              (terminated)
		);

	new_sdram_controller_grms_s1_translator : component p2_grms_qsys_new_sdram_controller_grms_s1_translator
		generic map (
			AV_ADDRESS_W                   => 22,
			AV_DATA_W                      => 16,
			UAV_DATA_W                     => 16,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 2,
			UAV_BYTEENABLE_W               => 2,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 2,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 1,
			USE_WAITREQUEST                => 1,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 2,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                                                 --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                          --                    reset.reset
			uav_address              => new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => new_sdram_controller_grms_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => new_sdram_controller_grms_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => new_sdram_controller_grms_s1_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => new_sdram_controller_grms_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => new_sdram_controller_grms_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_byteenable            => new_sdram_controller_grms_s1_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_readdatavalid         => new_sdram_controller_grms_s1_translator_avalon_anti_slave_0_readdatavalid,               --                         .readdatavalid
			av_waitrequest           => new_sdram_controller_grms_s1_translator_avalon_anti_slave_0_waitrequest,                 --                         .waitrequest
			av_chipselect            => new_sdram_controller_grms_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_begintransfer         => open,                                                                                    --              (terminated)
			av_beginbursttransfer    => open,                                                                                    --              (terminated)
			av_burstcount            => open,                                                                                    --              (terminated)
			av_writebyteenable       => open,                                                                                    --              (terminated)
			av_lock                  => open,                                                                                    --              (terminated)
			av_clken                 => open,                                                                                    --              (terminated)
			uav_clken                => '0',                                                                                     --              (terminated)
			av_debugaccess           => open,                                                                                    --              (terminated)
			av_outputenable          => open,                                                                                    --              (terminated)
			uav_response             => open,                                                                                    --              (terminated)
			av_response              => "00",                                                                                    --              (terminated)
			uav_writeresponserequest => '0',                                                                                     --              (terminated)
			uav_writeresponsevalid   => open,                                                                                    --              (terminated)
			av_writeresponserequest  => open,                                                                                    --              (terminated)
			av_writeresponsevalid    => '0'                                                                                      --              (terminated)
		);

	timer_grms_s1_translator : component p2_grms_qsys_timer_grms_s1_translator
		generic map (
			AV_ADDRESS_W                   => 3,
			AV_DATA_W                      => 16,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                                  --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                           --                    reset.reset
			uav_address              => timer_grms_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => timer_grms_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => timer_grms_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => timer_grms_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => timer_grms_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => timer_grms_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => timer_grms_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => timer_grms_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => timer_grms_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => timer_grms_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => timer_grms_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => timer_grms_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => timer_grms_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => timer_grms_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => timer_grms_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => timer_grms_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                     --              (terminated)
			av_begintransfer         => open,                                                                     --              (terminated)
			av_beginbursttransfer    => open,                                                                     --              (terminated)
			av_burstcount            => open,                                                                     --              (terminated)
			av_byteenable            => open,                                                                     --              (terminated)
			av_readdatavalid         => '0',                                                                      --              (terminated)
			av_waitrequest           => '0',                                                                      --              (terminated)
			av_writebyteenable       => open,                                                                     --              (terminated)
			av_lock                  => open,                                                                     --              (terminated)
			av_clken                 => open,                                                                     --              (terminated)
			uav_clken                => '0',                                                                      --              (terminated)
			av_debugaccess           => open,                                                                     --              (terminated)
			av_outputenable          => open,                                                                     --              (terminated)
			uav_response             => open,                                                                     --              (terminated)
			av_response              => "00",                                                                     --              (terminated)
			uav_writeresponserequest => '0',                                                                      --              (terminated)
			uav_writeresponsevalid   => open,                                                                     --              (terminated)
			av_writeresponserequest  => open,                                                                     --              (terminated)
			av_writeresponsevalid    => '0'                                                                       --              (terminated)
		);

	lcd_16207_grms_control_slave_translator : component p2_grms_qsys_lcd_16207_grms_control_slave_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 8,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 13,
			AV_WRITE_WAIT_CYCLES           => 13,
			AV_SETUP_WAIT_CYCLES           => 13,
			AV_DATA_HOLD_CYCLES            => 13
		)
		port map (
			clk                      => clk_clk,                                                                                 --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                          --                    reset.reset
			uav_address              => lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => lcd_16207_grms_control_slave_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => lcd_16207_grms_control_slave_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => lcd_16207_grms_control_slave_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => lcd_16207_grms_control_slave_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => lcd_16207_grms_control_slave_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_begintransfer         => lcd_16207_grms_control_slave_translator_avalon_anti_slave_0_begintransfer,               --                         .begintransfer
			av_beginbursttransfer    => open,                                                                                    --              (terminated)
			av_burstcount            => open,                                                                                    --              (terminated)
			av_byteenable            => open,                                                                                    --              (terminated)
			av_readdatavalid         => '0',                                                                                     --              (terminated)
			av_waitrequest           => '0',                                                                                     --              (terminated)
			av_writebyteenable       => open,                                                                                    --              (terminated)
			av_lock                  => open,                                                                                    --              (terminated)
			av_chipselect            => open,                                                                                    --              (terminated)
			av_clken                 => open,                                                                                    --              (terminated)
			uav_clken                => '0',                                                                                     --              (terminated)
			av_debugaccess           => open,                                                                                    --              (terminated)
			av_outputenable          => open,                                                                                    --              (terminated)
			uav_response             => open,                                                                                    --              (terminated)
			av_response              => "00",                                                                                    --              (terminated)
			uav_writeresponserequest => '0',                                                                                     --              (terminated)
			uav_writeresponsevalid   => open,                                                                                    --              (terminated)
			av_writeresponserequest  => open,                                                                                    --              (terminated)
			av_writeresponsevalid    => '0'                                                                                      --              (terminated)
		);

	pa_grms_s1_translator : component p2_grms_qsys_pa_grms_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                               --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                        --                    reset.reset
			uav_address              => pa_grms_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => pa_grms_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => pa_grms_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => pa_grms_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => pa_grms_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => pa_grms_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => pa_grms_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => pa_grms_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => pa_grms_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => pa_grms_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => pa_grms_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => pa_grms_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_readdata              => pa_grms_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_write                 => open,                                                                  --              (terminated)
			av_read                  => open,                                                                  --              (terminated)
			av_writedata             => open,                                                                  --              (terminated)
			av_begintransfer         => open,                                                                  --              (terminated)
			av_beginbursttransfer    => open,                                                                  --              (terminated)
			av_burstcount            => open,                                                                  --              (terminated)
			av_byteenable            => open,                                                                  --              (terminated)
			av_readdatavalid         => '0',                                                                   --              (terminated)
			av_waitrequest           => '0',                                                                   --              (terminated)
			av_writebyteenable       => open,                                                                  --              (terminated)
			av_lock                  => open,                                                                  --              (terminated)
			av_chipselect            => open,                                                                  --              (terminated)
			av_clken                 => open,                                                                  --              (terminated)
			uav_clken                => '0',                                                                   --              (terminated)
			av_debugaccess           => open,                                                                  --              (terminated)
			av_outputenable          => open,                                                                  --              (terminated)
			uav_response             => open,                                                                  --              (terminated)
			av_response              => "00",                                                                  --              (terminated)
			uav_writeresponserequest => '0',                                                                   --              (terminated)
			uav_writeresponsevalid   => open,                                                                  --              (terminated)
			av_writeresponserequest  => open,                                                                  --              (terminated)
			av_writeresponsevalid    => '0'                                                                    --              (terminated)
		);

	pb_grms_s1_translator : component p2_grms_qsys_pa_grms_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                               --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                        --                    reset.reset
			uav_address              => pb_grms_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => pb_grms_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => pb_grms_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => pb_grms_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => pb_grms_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => pb_grms_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => pb_grms_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => pb_grms_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => pb_grms_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => pb_grms_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => pb_grms_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => pb_grms_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_readdata              => pb_grms_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_write                 => open,                                                                  --              (terminated)
			av_read                  => open,                                                                  --              (terminated)
			av_writedata             => open,                                                                  --              (terminated)
			av_begintransfer         => open,                                                                  --              (terminated)
			av_beginbursttransfer    => open,                                                                  --              (terminated)
			av_burstcount            => open,                                                                  --              (terminated)
			av_byteenable            => open,                                                                  --              (terminated)
			av_readdatavalid         => '0',                                                                   --              (terminated)
			av_waitrequest           => '0',                                                                   --              (terminated)
			av_writebyteenable       => open,                                                                  --              (terminated)
			av_lock                  => open,                                                                  --              (terminated)
			av_chipselect            => open,                                                                  --              (terminated)
			av_clken                 => open,                                                                  --              (terminated)
			uav_clken                => '0',                                                                   --              (terminated)
			av_debugaccess           => open,                                                                  --              (terminated)
			av_outputenable          => open,                                                                  --              (terminated)
			uav_response             => open,                                                                  --              (terminated)
			av_response              => "00",                                                                  --              (terminated)
			uav_writeresponserequest => '0',                                                                   --              (terminated)
			uav_writeresponsevalid   => open,                                                                  --              (terminated)
			av_writeresponserequest  => open,                                                                  --              (terminated)
			av_writeresponsevalid    => '0'                                                                    --              (terminated)
		);

	pc_grms_s1_translator : component p2_grms_qsys_pc_grms_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                               --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                        --                    reset.reset
			uav_address              => pc_grms_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => pc_grms_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => pc_grms_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => pc_grms_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => pc_grms_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => pc_grms_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => pc_grms_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => pc_grms_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => pc_grms_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => pc_grms_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => pc_grms_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => pc_grms_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => pc_grms_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => pc_grms_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => pc_grms_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => pc_grms_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                  --              (terminated)
			av_begintransfer         => open,                                                                  --              (terminated)
			av_beginbursttransfer    => open,                                                                  --              (terminated)
			av_burstcount            => open,                                                                  --              (terminated)
			av_byteenable            => open,                                                                  --              (terminated)
			av_readdatavalid         => '0',                                                                   --              (terminated)
			av_waitrequest           => '0',                                                                   --              (terminated)
			av_writebyteenable       => open,                                                                  --              (terminated)
			av_lock                  => open,                                                                  --              (terminated)
			av_clken                 => open,                                                                  --              (terminated)
			uav_clken                => '0',                                                                   --              (terminated)
			av_debugaccess           => open,                                                                  --              (terminated)
			av_outputenable          => open,                                                                  --              (terminated)
			uav_response             => open,                                                                  --              (terminated)
			av_response              => "00",                                                                  --              (terminated)
			uav_writeresponserequest => '0',                                                                   --              (terminated)
			uav_writeresponsevalid   => open,                                                                  --              (terminated)
			av_writeresponserequest  => open,                                                                  --              (terminated)
			av_writeresponsevalid    => '0'                                                                    --              (terminated)
		);

	pd_grms_s1_translator : component p2_grms_qsys_pc_grms_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                               --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                        --                    reset.reset
			uav_address              => pd_grms_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => pd_grms_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => pd_grms_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => pd_grms_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => pd_grms_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => pd_grms_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => pd_grms_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => pd_grms_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => pd_grms_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => pd_grms_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => pd_grms_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => pd_grms_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => pd_grms_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => pd_grms_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => pd_grms_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => pd_grms_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                  --              (terminated)
			av_begintransfer         => open,                                                                  --              (terminated)
			av_beginbursttransfer    => open,                                                                  --              (terminated)
			av_burstcount            => open,                                                                  --              (terminated)
			av_byteenable            => open,                                                                  --              (terminated)
			av_readdatavalid         => '0',                                                                   --              (terminated)
			av_waitrequest           => '0',                                                                   --              (terminated)
			av_writebyteenable       => open,                                                                  --              (terminated)
			av_lock                  => open,                                                                  --              (terminated)
			av_clken                 => open,                                                                  --              (terminated)
			uav_clken                => '0',                                                                   --              (terminated)
			av_debugaccess           => open,                                                                  --              (terminated)
			av_outputenable          => open,                                                                  --              (terminated)
			uav_response             => open,                                                                  --              (terminated)
			av_response              => "00",                                                                  --              (terminated)
			uav_writeresponserequest => '0',                                                                   --              (terminated)
			uav_writeresponsevalid   => open,                                                                  --              (terminated)
			av_writeresponserequest  => open,                                                                  --              (terminated)
			av_writeresponsevalid    => '0'                                                                    --              (terminated)
		);

	pe_grms_s1_translator : component p2_grms_qsys_pc_grms_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                               --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                        --                    reset.reset
			uav_address              => pe_grms_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => pe_grms_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => pe_grms_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => pe_grms_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => pe_grms_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => pe_grms_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => pe_grms_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => pe_grms_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => pe_grms_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => pe_grms_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => pe_grms_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => pe_grms_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => pe_grms_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => pe_grms_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => pe_grms_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => pe_grms_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                  --              (terminated)
			av_begintransfer         => open,                                                                  --              (terminated)
			av_beginbursttransfer    => open,                                                                  --              (terminated)
			av_burstcount            => open,                                                                  --              (terminated)
			av_byteenable            => open,                                                                  --              (terminated)
			av_readdatavalid         => '0',                                                                   --              (terminated)
			av_waitrequest           => '0',                                                                   --              (terminated)
			av_writebyteenable       => open,                                                                  --              (terminated)
			av_lock                  => open,                                                                  --              (terminated)
			av_clken                 => open,                                                                  --              (terminated)
			uav_clken                => '0',                                                                   --              (terminated)
			av_debugaccess           => open,                                                                  --              (terminated)
			av_outputenable          => open,                                                                  --              (terminated)
			uav_response             => open,                                                                  --              (terminated)
			av_response              => "00",                                                                  --              (terminated)
			uav_writeresponserequest => '0',                                                                   --              (terminated)
			uav_writeresponsevalid   => open,                                                                  --              (terminated)
			av_writeresponserequest  => open,                                                                  --              (terminated)
			av_writeresponsevalid    => '0'                                                                    --              (terminated)
		);

	pf_grms_s1_translator : component p2_grms_qsys_pc_grms_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                               --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                        --                    reset.reset
			uav_address              => pf_grms_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => pf_grms_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => pf_grms_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => pf_grms_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => pf_grms_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => pf_grms_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => pf_grms_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => pf_grms_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => pf_grms_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => pf_grms_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => pf_grms_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => pf_grms_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => pf_grms_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => pf_grms_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => pf_grms_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => pf_grms_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                  --              (terminated)
			av_begintransfer         => open,                                                                  --              (terminated)
			av_beginbursttransfer    => open,                                                                  --              (terminated)
			av_burstcount            => open,                                                                  --              (terminated)
			av_byteenable            => open,                                                                  --              (terminated)
			av_readdatavalid         => '0',                                                                   --              (terminated)
			av_waitrequest           => '0',                                                                   --              (terminated)
			av_writebyteenable       => open,                                                                  --              (terminated)
			av_lock                  => open,                                                                  --              (terminated)
			av_clken                 => open,                                                                  --              (terminated)
			uav_clken                => '0',                                                                   --              (terminated)
			av_debugaccess           => open,                                                                  --              (terminated)
			av_outputenable          => open,                                                                  --              (terminated)
			uav_response             => open,                                                                  --              (terminated)
			av_response              => "00",                                                                  --              (terminated)
			uav_writeresponserequest => '0',                                                                   --              (terminated)
			uav_writeresponsevalid   => open,                                                                  --              (terminated)
			av_writeresponserequest  => open,                                                                  --              (terminated)
			av_writeresponsevalid    => '0'                                                                    --              (terminated)
		);

	pg_grms_s1_translator : component p2_grms_qsys_pc_grms_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                               --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                        --                    reset.reset
			uav_address              => pg_grms_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => pg_grms_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => pg_grms_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => pg_grms_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => pg_grms_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => pg_grms_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => pg_grms_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => pg_grms_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => pg_grms_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => pg_grms_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => pg_grms_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => pg_grms_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => pg_grms_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => pg_grms_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => pg_grms_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => pg_grms_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                  --              (terminated)
			av_begintransfer         => open,                                                                  --              (terminated)
			av_beginbursttransfer    => open,                                                                  --              (terminated)
			av_burstcount            => open,                                                                  --              (terminated)
			av_byteenable            => open,                                                                  --              (terminated)
			av_readdatavalid         => '0',                                                                   --              (terminated)
			av_waitrequest           => '0',                                                                   --              (terminated)
			av_writebyteenable       => open,                                                                  --              (terminated)
			av_lock                  => open,                                                                  --              (terminated)
			av_clken                 => open,                                                                  --              (terminated)
			uav_clken                => '0',                                                                   --              (terminated)
			av_debugaccess           => open,                                                                  --              (terminated)
			av_outputenable          => open,                                                                  --              (terminated)
			uav_response             => open,                                                                  --              (terminated)
			av_response              => "00",                                                                  --              (terminated)
			uav_writeresponserequest => '0',                                                                   --              (terminated)
			uav_writeresponsevalid   => open,                                                                  --              (terminated)
			av_writeresponserequest  => open,                                                                  --              (terminated)
			av_writeresponsevalid    => '0'                                                                    --              (terminated)
		);

	ph_grms_s1_translator : component p2_grms_qsys_pc_grms_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                               --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                        --                    reset.reset
			uav_address              => ph_grms_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => ph_grms_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => ph_grms_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => ph_grms_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => ph_grms_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => ph_grms_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => ph_grms_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => ph_grms_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => ph_grms_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => ph_grms_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => ph_grms_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => ph_grms_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => ph_grms_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => ph_grms_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => ph_grms_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => ph_grms_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                  --              (terminated)
			av_begintransfer         => open,                                                                  --              (terminated)
			av_beginbursttransfer    => open,                                                                  --              (terminated)
			av_burstcount            => open,                                                                  --              (terminated)
			av_byteenable            => open,                                                                  --              (terminated)
			av_readdatavalid         => '0',                                                                   --              (terminated)
			av_waitrequest           => '0',                                                                   --              (terminated)
			av_writebyteenable       => open,                                                                  --              (terminated)
			av_lock                  => open,                                                                  --              (terminated)
			av_clken                 => open,                                                                  --              (terminated)
			uav_clken                => '0',                                                                   --              (terminated)
			av_debugaccess           => open,                                                                  --              (terminated)
			av_outputenable          => open,                                                                  --              (terminated)
			uav_response             => open,                                                                  --              (terminated)
			av_response              => "00",                                                                  --              (terminated)
			uav_writeresponserequest => '0',                                                                   --              (terminated)
			uav_writeresponsevalid   => open,                                                                  --              (terminated)
			av_writeresponserequest  => open,                                                                  --              (terminated)
			av_writeresponsevalid    => '0'                                                                    --              (terminated)
		);

	pi_grms_s1_translator : component p2_grms_qsys_pc_grms_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                               --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                        --                    reset.reset
			uav_address              => pi_grms_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => pi_grms_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => pi_grms_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => pi_grms_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => pi_grms_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => pi_grms_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => pi_grms_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => pi_grms_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => pi_grms_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => pi_grms_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => pi_grms_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => pi_grms_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => pi_grms_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => pi_grms_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => pi_grms_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => pi_grms_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                  --              (terminated)
			av_begintransfer         => open,                                                                  --              (terminated)
			av_beginbursttransfer    => open,                                                                  --              (terminated)
			av_burstcount            => open,                                                                  --              (terminated)
			av_byteenable            => open,                                                                  --              (terminated)
			av_readdatavalid         => '0',                                                                   --              (terminated)
			av_waitrequest           => '0',                                                                   --              (terminated)
			av_writebyteenable       => open,                                                                  --              (terminated)
			av_lock                  => open,                                                                  --              (terminated)
			av_clken                 => open,                                                                  --              (terminated)
			uav_clken                => '0',                                                                   --              (terminated)
			av_debugaccess           => open,                                                                  --              (terminated)
			av_outputenable          => open,                                                                  --              (terminated)
			uav_response             => open,                                                                  --              (terminated)
			av_response              => "00",                                                                  --              (terminated)
			uav_writeresponserequest => '0',                                                                   --              (terminated)
			uav_writeresponsevalid   => open,                                                                  --              (terminated)
			av_writeresponserequest  => open,                                                                  --              (terminated)
			av_writeresponsevalid    => '0'                                                                    --              (terminated)
		);

	nios2_qsys_grms_instruction_master_translator_avalon_universal_master_0_agent : component altera_merlin_master_agent
		generic map (
			PKT_PROTECTION_H          => 93,
			PKT_PROTECTION_L          => 91,
			PKT_BEGIN_BURST           => 80,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			PKT_BURST_TYPE_H          => 77,
			PKT_BURST_TYPE_L          => 76,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_TRANS_EXCLUSIVE       => 66,
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_SRC_ID_H              => 85,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 89,
			PKT_DEST_ID_L             => 86,
			PKT_THREAD_ID_H           => 90,
			PKT_THREAD_ID_L           => 90,
			PKT_CACHE_H               => 97,
			PKT_CACHE_L               => 94,
			PKT_DATA_SIDEBAND_H       => 79,
			PKT_DATA_SIDEBAND_L       => 79,
			PKT_QOS_H                 => 81,
			PKT_QOS_L                 => 81,
			PKT_ADDR_SIDEBAND_H       => 78,
			PKT_ADDR_SIDEBAND_L       => 78,
			PKT_RESPONSE_STATUS_H     => 99,
			PKT_RESPONSE_STATUS_L     => 98,
			ST_DATA_W                 => 100,
			ST_CHANNEL_W              => 14,
			AV_BURSTCOUNT_W           => 3,
			SUPPRESS_0_BYTEEN_RSP     => 0,
			ID                        => 1,
			BURSTWRAP_VALUE           => 3,
			CACHE_VALUE               => 0,
			SECURE_ACCESS_BIT         => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                                        --       clk.clk
			reset                   => rst_controller_reset_out_reset,                                                                 -- clk_reset.reset
			av_address              => nios2_qsys_grms_instruction_master_translator_avalon_universal_master_0_address,                --        av.address
			av_write                => nios2_qsys_grms_instruction_master_translator_avalon_universal_master_0_write,                  --          .write
			av_read                 => nios2_qsys_grms_instruction_master_translator_avalon_universal_master_0_read,                   --          .read
			av_writedata            => nios2_qsys_grms_instruction_master_translator_avalon_universal_master_0_writedata,              --          .writedata
			av_readdata             => nios2_qsys_grms_instruction_master_translator_avalon_universal_master_0_readdata,               --          .readdata
			av_waitrequest          => nios2_qsys_grms_instruction_master_translator_avalon_universal_master_0_waitrequest,            --          .waitrequest
			av_readdatavalid        => nios2_qsys_grms_instruction_master_translator_avalon_universal_master_0_readdatavalid,          --          .readdatavalid
			av_byteenable           => nios2_qsys_grms_instruction_master_translator_avalon_universal_master_0_byteenable,             --          .byteenable
			av_burstcount           => nios2_qsys_grms_instruction_master_translator_avalon_universal_master_0_burstcount,             --          .burstcount
			av_debugaccess          => nios2_qsys_grms_instruction_master_translator_avalon_universal_master_0_debugaccess,            --          .debugaccess
			av_lock                 => nios2_qsys_grms_instruction_master_translator_avalon_universal_master_0_lock,                   --          .lock
			cp_valid                => nios2_qsys_grms_instruction_master_translator_avalon_universal_master_0_agent_cp_valid,         --        cp.valid
			cp_data                 => nios2_qsys_grms_instruction_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			cp_startofpacket        => nios2_qsys_grms_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			cp_endofpacket          => nios2_qsys_grms_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			cp_ready                => nios2_qsys_grms_instruction_master_translator_avalon_universal_master_0_agent_cp_ready,         --          .ready
			rp_valid                => rsp_xbar_mux_src_valid,                                                                         --        rp.valid
			rp_data                 => rsp_xbar_mux_src_data,                                                                          --          .data
			rp_channel              => rsp_xbar_mux_src_channel,                                                                       --          .channel
			rp_startofpacket        => rsp_xbar_mux_src_startofpacket,                                                                 --          .startofpacket
			rp_endofpacket          => rsp_xbar_mux_src_endofpacket,                                                                   --          .endofpacket
			rp_ready                => rsp_xbar_mux_src_ready,                                                                         --          .ready
			av_response             => open,                                                                                           -- (terminated)
			av_writeresponserequest => '0',                                                                                            -- (terminated)
			av_writeresponsevalid   => open                                                                                            -- (terminated)
		);

	nios2_qsys_grms_data_master_translator_avalon_universal_master_0_agent : component altera_merlin_master_agent
		generic map (
			PKT_PROTECTION_H          => 93,
			PKT_PROTECTION_L          => 91,
			PKT_BEGIN_BURST           => 80,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			PKT_BURST_TYPE_H          => 77,
			PKT_BURST_TYPE_L          => 76,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_TRANS_EXCLUSIVE       => 66,
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_SRC_ID_H              => 85,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 89,
			PKT_DEST_ID_L             => 86,
			PKT_THREAD_ID_H           => 90,
			PKT_THREAD_ID_L           => 90,
			PKT_CACHE_H               => 97,
			PKT_CACHE_L               => 94,
			PKT_DATA_SIDEBAND_H       => 79,
			PKT_DATA_SIDEBAND_L       => 79,
			PKT_QOS_H                 => 81,
			PKT_QOS_L                 => 81,
			PKT_ADDR_SIDEBAND_H       => 78,
			PKT_ADDR_SIDEBAND_L       => 78,
			PKT_RESPONSE_STATUS_H     => 99,
			PKT_RESPONSE_STATUS_L     => 98,
			ST_DATA_W                 => 100,
			ST_CHANNEL_W              => 14,
			AV_BURSTCOUNT_W           => 3,
			SUPPRESS_0_BYTEEN_RSP     => 0,
			ID                        => 0,
			BURSTWRAP_VALUE           => 7,
			CACHE_VALUE               => 0,
			SECURE_ACCESS_BIT         => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                                 --       clk.clk
			reset                   => rst_controller_reset_out_reset,                                                          -- clk_reset.reset
			av_address              => nios2_qsys_grms_data_master_translator_avalon_universal_master_0_address,                --        av.address
			av_write                => nios2_qsys_grms_data_master_translator_avalon_universal_master_0_write,                  --          .write
			av_read                 => nios2_qsys_grms_data_master_translator_avalon_universal_master_0_read,                   --          .read
			av_writedata            => nios2_qsys_grms_data_master_translator_avalon_universal_master_0_writedata,              --          .writedata
			av_readdata             => nios2_qsys_grms_data_master_translator_avalon_universal_master_0_readdata,               --          .readdata
			av_waitrequest          => nios2_qsys_grms_data_master_translator_avalon_universal_master_0_waitrequest,            --          .waitrequest
			av_readdatavalid        => nios2_qsys_grms_data_master_translator_avalon_universal_master_0_readdatavalid,          --          .readdatavalid
			av_byteenable           => nios2_qsys_grms_data_master_translator_avalon_universal_master_0_byteenable,             --          .byteenable
			av_burstcount           => nios2_qsys_grms_data_master_translator_avalon_universal_master_0_burstcount,             --          .burstcount
			av_debugaccess          => nios2_qsys_grms_data_master_translator_avalon_universal_master_0_debugaccess,            --          .debugaccess
			av_lock                 => nios2_qsys_grms_data_master_translator_avalon_universal_master_0_lock,                   --          .lock
			cp_valid                => nios2_qsys_grms_data_master_translator_avalon_universal_master_0_agent_cp_valid,         --        cp.valid
			cp_data                 => nios2_qsys_grms_data_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			cp_startofpacket        => nios2_qsys_grms_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			cp_endofpacket          => nios2_qsys_grms_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			cp_ready                => nios2_qsys_grms_data_master_translator_avalon_universal_master_0_agent_cp_ready,         --          .ready
			rp_valid                => rsp_xbar_mux_001_src_valid,                                                              --        rp.valid
			rp_data                 => rsp_xbar_mux_001_src_data,                                                               --          .data
			rp_channel              => rsp_xbar_mux_001_src_channel,                                                            --          .channel
			rp_startofpacket        => rsp_xbar_mux_001_src_startofpacket,                                                      --          .startofpacket
			rp_endofpacket          => rsp_xbar_mux_001_src_endofpacket,                                                        --          .endofpacket
			rp_ready                => rsp_xbar_mux_001_src_ready,                                                              --          .ready
			av_response             => open,                                                                                    -- (terminated)
			av_writeresponserequest => '0',                                                                                     -- (terminated)
			av_writeresponsevalid   => open                                                                                     -- (terminated)
		);

	nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent : component p2_grms_qsys_nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 85,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 89,
			PKT_DEST_ID_L             => 86,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 93,
			PKT_PROTECTION_L          => 91,
			PKT_RESPONSE_STATUS_H     => 99,
			PKT_RESPONSE_STATUS_L     => 98,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 14,
			ST_DATA_W                 => 100,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                                                --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                                         --       clk_reset.reset
			m0_address              => nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_src_ready,                                                                                 --              cp.ready
			cp_valid                => cmd_xbar_mux_src_valid,                                                                                 --                .valid
			cp_data                 => cmd_xbar_mux_src_data,                                                                                  --                .data
			cp_startofpacket        => cmd_xbar_mux_src_startofpacket,                                                                         --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_src_endofpacket,                                                                           --                .endofpacket
			cp_channel              => cmd_xbar_mux_src_channel,                                                                               --                .channel
			rf_sink_ready           => nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                                   --     (terminated)
			m0_writeresponserequest => open,                                                                                                   --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                                     --     (terminated)
		);

	nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo : component p2_grms_qsys_nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 101,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                                                --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                                         -- clk_reset.reset
			in_data           => nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                                   -- (terminated)
			csr_read          => '0',                                                                                                    -- (terminated)
			csr_write         => '0',                                                                                                    -- (terminated)
			csr_readdata      => open,                                                                                                   -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                                     -- (terminated)
			almost_full_data  => open,                                                                                                   -- (terminated)
			almost_empty_data => open,                                                                                                   -- (terminated)
			in_empty          => '0',                                                                                                    -- (terminated)
			out_empty         => open,                                                                                                   -- (terminated)
			in_error          => '0',                                                                                                    -- (terminated)
			out_error         => open,                                                                                                   -- (terminated)
			in_channel        => '0',                                                                                                    -- (terminated)
			out_channel       => open                                                                                                    -- (terminated)
		);

	jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent : component p2_grms_qsys_nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 85,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 89,
			PKT_DEST_ID_L             => 86,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 93,
			PKT_PROTECTION_L          => 91,
			PKT_RESPONSE_STATUS_H     => 99,
			PKT_RESPONSE_STATUS_L     => 98,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 14,
			ST_DATA_W                 => 100,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                                               --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                                        --       clk_reset.reset
			m0_address              => jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_001_src_ready,                                                                            --              cp.ready
			cp_valid                => cmd_xbar_mux_001_src_valid,                                                                            --                .valid
			cp_data                 => cmd_xbar_mux_001_src_data,                                                                             --                .data
			cp_startofpacket        => cmd_xbar_mux_001_src_startofpacket,                                                                    --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_001_src_endofpacket,                                                                      --                .endofpacket
			cp_channel              => cmd_xbar_mux_001_src_channel,                                                                          --                .channel
			rf_sink_ready           => jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                                  --     (terminated)
			m0_writeresponserequest => open,                                                                                                  --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                                    --     (terminated)
		);

	jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo : component p2_grms_qsys_nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 101,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                                               --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                                        -- clk_reset.reset
			in_data           => jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                                  -- (terminated)
			csr_read          => '0',                                                                                                   -- (terminated)
			csr_write         => '0',                                                                                                   -- (terminated)
			csr_readdata      => open,                                                                                                  -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                                    -- (terminated)
			almost_full_data  => open,                                                                                                  -- (terminated)
			almost_empty_data => open,                                                                                                  -- (terminated)
			in_empty          => '0',                                                                                                   -- (terminated)
			out_empty         => open,                                                                                                  -- (terminated)
			in_error          => '0',                                                                                                   -- (terminated)
			out_error         => open,                                                                                                  -- (terminated)
			in_channel        => '0',                                                                                                   -- (terminated)
			out_channel       => open                                                                                                   -- (terminated)
		);

	new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent : component p2_grms_qsys_new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 15,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 62,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 17,
			PKT_BYTEEN_L              => 16,
			PKT_ADDR_H                => 42,
			PKT_ADDR_L                => 18,
			PKT_TRANS_COMPRESSED_READ => 43,
			PKT_TRANS_POSTED          => 44,
			PKT_TRANS_WRITE           => 45,
			PKT_TRANS_READ            => 46,
			PKT_TRANS_LOCK            => 47,
			PKT_SRC_ID_H              => 67,
			PKT_SRC_ID_L              => 64,
			PKT_DEST_ID_H             => 71,
			PKT_DEST_ID_L             => 68,
			PKT_BURSTWRAP_H           => 54,
			PKT_BURSTWRAP_L           => 52,
			PKT_BYTE_CNT_H            => 51,
			PKT_BYTE_CNT_L            => 49,
			PKT_PROTECTION_H          => 75,
			PKT_PROTECTION_L          => 73,
			PKT_RESPONSE_STATUS_H     => 81,
			PKT_RESPONSE_STATUS_L     => 80,
			PKT_BURST_SIZE_H          => 57,
			PKT_BURST_SIZE_L          => 55,
			ST_CHANNEL_W              => 14,
			ST_DATA_W                 => 82,
			AVS_BURSTCOUNT_W          => 2,
			SUPPRESS_0_BYTEEN_CMD     => 1,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                                           --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                                    --       clk_reset.reset
			m0_address              => new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => burst_adapter_source0_ready,                                                                       --              cp.ready
			cp_valid                => burst_adapter_source0_valid,                                                                       --                .valid
			cp_data                 => burst_adapter_source0_data,                                                                        --                .data
			cp_startofpacket        => burst_adapter_source0_startofpacket,                                                               --                .startofpacket
			cp_endofpacket          => burst_adapter_source0_endofpacket,                                                                 --                .endofpacket
			cp_channel              => burst_adapter_source0_channel,                                                                     --                .channel
			rf_sink_ready           => new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid,       --                .valid
			rdata_fifo_sink_data    => new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,        --                .data
			rdata_fifo_src_ready    => new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                              --     (terminated)
			m0_writeresponserequest => open,                                                                                              --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                                --     (terminated)
		);

	new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component p2_grms_qsys_new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 83,
			FIFO_DEPTH          => 8,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                                           --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                                    -- clk_reset.reset
			in_data           => new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                              -- (terminated)
			csr_read          => '0',                                                                                               -- (terminated)
			csr_write         => '0',                                                                                               -- (terminated)
			csr_readdata      => open,                                                                                              -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                                -- (terminated)
			almost_full_data  => open,                                                                                              -- (terminated)
			almost_empty_data => open,                                                                                              -- (terminated)
			in_empty          => '0',                                                                                               -- (terminated)
			out_empty         => open,                                                                                              -- (terminated)
			in_error          => '0',                                                                                               -- (terminated)
			out_error         => open,                                                                                              -- (terminated)
			in_channel        => '0',                                                                                               -- (terminated)
			out_channel       => open                                                                                               -- (terminated)
		);

	new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo : component p2_grms_qsys_new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 18,
			FIFO_DEPTH          => 8,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 0,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 3,
			USE_MEMORY_BLOCKS   => 1,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                                     --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                              -- clk_reset.reset
			in_data           => new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,  --        in.data
			in_valid          => new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid, --          .valid
			in_ready          => new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready, --          .ready
			out_data          => new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,  --       out.data
			out_valid         => new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid, --          .valid
			out_ready         => new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready, --          .ready
			csr_address       => "00",                                                                                        -- (terminated)
			csr_read          => '0',                                                                                         -- (terminated)
			csr_write         => '0',                                                                                         -- (terminated)
			csr_readdata      => open,                                                                                        -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                          -- (terminated)
			almost_full_data  => open,                                                                                        -- (terminated)
			almost_empty_data => open,                                                                                        -- (terminated)
			in_startofpacket  => '0',                                                                                         -- (terminated)
			in_endofpacket    => '0',                                                                                         -- (terminated)
			out_startofpacket => open,                                                                                        -- (terminated)
			out_endofpacket   => open,                                                                                        -- (terminated)
			in_empty          => '0',                                                                                         -- (terminated)
			out_empty         => open,                                                                                        -- (terminated)
			in_error          => '0',                                                                                         -- (terminated)
			out_error         => open,                                                                                        -- (terminated)
			in_channel        => '0',                                                                                         -- (terminated)
			out_channel       => open                                                                                         -- (terminated)
		);

	timer_grms_s1_translator_avalon_universal_slave_0_agent : component p2_grms_qsys_nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 85,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 89,
			PKT_DEST_ID_L             => 86,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 93,
			PKT_PROTECTION_L          => 91,
			PKT_RESPONSE_STATUS_H     => 99,
			PKT_RESPONSE_STATUS_L     => 98,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 14,
			ST_DATA_W                 => 100,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                            --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                     --       clk_reset.reset
			m0_address              => timer_grms_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => timer_grms_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => timer_grms_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => timer_grms_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => timer_grms_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => timer_grms_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => timer_grms_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => timer_grms_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => timer_grms_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => timer_grms_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => timer_grms_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => timer_grms_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => timer_grms_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => timer_grms_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => timer_grms_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => timer_grms_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_003_src_ready,                                                         --              cp.ready
			cp_valid                => cmd_xbar_mux_003_src_valid,                                                         --                .valid
			cp_data                 => cmd_xbar_mux_003_src_data,                                                          --                .data
			cp_startofpacket        => cmd_xbar_mux_003_src_startofpacket,                                                 --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_003_src_endofpacket,                                                   --                .endofpacket
			cp_channel              => cmd_xbar_mux_003_src_channel,                                                       --                .channel
			rf_sink_ready           => timer_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => timer_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => timer_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => timer_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => timer_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => timer_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => timer_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => timer_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => timer_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => timer_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => timer_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => timer_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => timer_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => timer_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => timer_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => timer_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                               --     (terminated)
			m0_writeresponserequest => open,                                                                               --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                 --     (terminated)
		);

	timer_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component p2_grms_qsys_nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 101,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                            --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                     -- clk_reset.reset
			in_data           => timer_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => timer_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => timer_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => timer_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => timer_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => timer_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => timer_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => timer_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => timer_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => timer_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                               -- (terminated)
			csr_read          => '0',                                                                                -- (terminated)
			csr_write         => '0',                                                                                -- (terminated)
			csr_readdata      => open,                                                                               -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                 -- (terminated)
			almost_full_data  => open,                                                                               -- (terminated)
			almost_empty_data => open,                                                                               -- (terminated)
			in_empty          => '0',                                                                                -- (terminated)
			out_empty         => open,                                                                               -- (terminated)
			in_error          => '0',                                                                                -- (terminated)
			out_error         => open,                                                                               -- (terminated)
			in_channel        => '0',                                                                                -- (terminated)
			out_channel       => open                                                                                -- (terminated)
		);

	lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent : component p2_grms_qsys_nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 85,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 89,
			PKT_DEST_ID_L             => 86,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 93,
			PKT_PROTECTION_L          => 91,
			PKT_RESPONSE_STATUS_H     => 99,
			PKT_RESPONSE_STATUS_L     => 98,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 14,
			ST_DATA_W                 => 100,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                                           --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                                    --       clk_reset.reset
			m0_address              => lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_004_src_ready,                                                                        --              cp.ready
			cp_valid                => cmd_xbar_mux_004_src_valid,                                                                        --                .valid
			cp_data                 => cmd_xbar_mux_004_src_data,                                                                         --                .data
			cp_startofpacket        => cmd_xbar_mux_004_src_startofpacket,                                                                --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_004_src_endofpacket,                                                                  --                .endofpacket
			cp_channel              => cmd_xbar_mux_004_src_channel,                                                                      --                .channel
			rf_sink_ready           => lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                              --     (terminated)
			m0_writeresponserequest => open,                                                                                              --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                                --     (terminated)
		);

	lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo : component p2_grms_qsys_nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 101,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                                           --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                                    -- clk_reset.reset
			in_data           => lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                              -- (terminated)
			csr_read          => '0',                                                                                               -- (terminated)
			csr_write         => '0',                                                                                               -- (terminated)
			csr_readdata      => open,                                                                                              -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                                -- (terminated)
			almost_full_data  => open,                                                                                              -- (terminated)
			almost_empty_data => open,                                                                                              -- (terminated)
			in_empty          => '0',                                                                                               -- (terminated)
			out_empty         => open,                                                                                              -- (terminated)
			in_error          => '0',                                                                                               -- (terminated)
			out_error         => open,                                                                                              -- (terminated)
			in_channel        => '0',                                                                                               -- (terminated)
			out_channel       => open                                                                                               -- (terminated)
		);

	pa_grms_s1_translator_avalon_universal_slave_0_agent : component p2_grms_qsys_nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 85,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 89,
			PKT_DEST_ID_L             => 86,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 93,
			PKT_PROTECTION_L          => 91,
			PKT_RESPONSE_STATUS_H     => 99,
			PKT_RESPONSE_STATUS_L     => 98,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 14,
			ST_DATA_W                 => 100,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                         --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                  --       clk_reset.reset
			m0_address              => pa_grms_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => pa_grms_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => pa_grms_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => pa_grms_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => pa_grms_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => pa_grms_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => pa_grms_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => pa_grms_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => pa_grms_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => pa_grms_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => pa_grms_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => pa_grms_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => pa_grms_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => pa_grms_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => pa_grms_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => pa_grms_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_005_src_ready,                                                      --              cp.ready
			cp_valid                => cmd_xbar_mux_005_src_valid,                                                      --                .valid
			cp_data                 => cmd_xbar_mux_005_src_data,                                                       --                .data
			cp_startofpacket        => cmd_xbar_mux_005_src_startofpacket,                                              --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_005_src_endofpacket,                                                --                .endofpacket
			cp_channel              => cmd_xbar_mux_005_src_channel,                                                    --                .channel
			rf_sink_ready           => pa_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => pa_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => pa_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => pa_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => pa_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => pa_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => pa_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => pa_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => pa_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => pa_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => pa_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => pa_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => pa_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => pa_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => pa_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => pa_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                            --     (terminated)
			m0_writeresponserequest => open,                                                                            --     (terminated)
			m0_writeresponsevalid   => '0'                                                                              --     (terminated)
		);

	pa_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component p2_grms_qsys_nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 101,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                         --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                  -- clk_reset.reset
			in_data           => pa_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => pa_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => pa_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => pa_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => pa_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => pa_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => pa_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => pa_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => pa_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => pa_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                            -- (terminated)
			csr_read          => '0',                                                                             -- (terminated)
			csr_write         => '0',                                                                             -- (terminated)
			csr_readdata      => open,                                                                            -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                              -- (terminated)
			almost_full_data  => open,                                                                            -- (terminated)
			almost_empty_data => open,                                                                            -- (terminated)
			in_empty          => '0',                                                                             -- (terminated)
			out_empty         => open,                                                                            -- (terminated)
			in_error          => '0',                                                                             -- (terminated)
			out_error         => open,                                                                            -- (terminated)
			in_channel        => '0',                                                                             -- (terminated)
			out_channel       => open                                                                             -- (terminated)
		);

	pb_grms_s1_translator_avalon_universal_slave_0_agent : component p2_grms_qsys_nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 85,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 89,
			PKT_DEST_ID_L             => 86,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 93,
			PKT_PROTECTION_L          => 91,
			PKT_RESPONSE_STATUS_H     => 99,
			PKT_RESPONSE_STATUS_L     => 98,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 14,
			ST_DATA_W                 => 100,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                         --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                  --       clk_reset.reset
			m0_address              => pb_grms_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => pb_grms_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => pb_grms_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => pb_grms_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => pb_grms_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => pb_grms_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => pb_grms_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => pb_grms_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => pb_grms_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => pb_grms_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => pb_grms_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => pb_grms_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => pb_grms_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => pb_grms_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => pb_grms_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => pb_grms_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_006_src_ready,                                                      --              cp.ready
			cp_valid                => cmd_xbar_mux_006_src_valid,                                                      --                .valid
			cp_data                 => cmd_xbar_mux_006_src_data,                                                       --                .data
			cp_startofpacket        => cmd_xbar_mux_006_src_startofpacket,                                              --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_006_src_endofpacket,                                                --                .endofpacket
			cp_channel              => cmd_xbar_mux_006_src_channel,                                                    --                .channel
			rf_sink_ready           => pb_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => pb_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => pb_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => pb_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => pb_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => pb_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => pb_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => pb_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => pb_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => pb_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => pb_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => pb_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => pb_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => pb_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => pb_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => pb_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                            --     (terminated)
			m0_writeresponserequest => open,                                                                            --     (terminated)
			m0_writeresponsevalid   => '0'                                                                              --     (terminated)
		);

	pb_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component p2_grms_qsys_nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 101,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                         --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                  -- clk_reset.reset
			in_data           => pb_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => pb_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => pb_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => pb_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => pb_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => pb_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => pb_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => pb_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => pb_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => pb_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                            -- (terminated)
			csr_read          => '0',                                                                             -- (terminated)
			csr_write         => '0',                                                                             -- (terminated)
			csr_readdata      => open,                                                                            -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                              -- (terminated)
			almost_full_data  => open,                                                                            -- (terminated)
			almost_empty_data => open,                                                                            -- (terminated)
			in_empty          => '0',                                                                             -- (terminated)
			out_empty         => open,                                                                            -- (terminated)
			in_error          => '0',                                                                             -- (terminated)
			out_error         => open,                                                                            -- (terminated)
			in_channel        => '0',                                                                             -- (terminated)
			out_channel       => open                                                                             -- (terminated)
		);

	pc_grms_s1_translator_avalon_universal_slave_0_agent : component p2_grms_qsys_nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 85,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 89,
			PKT_DEST_ID_L             => 86,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 93,
			PKT_PROTECTION_L          => 91,
			PKT_RESPONSE_STATUS_H     => 99,
			PKT_RESPONSE_STATUS_L     => 98,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 14,
			ST_DATA_W                 => 100,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                         --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                  --       clk_reset.reset
			m0_address              => pc_grms_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => pc_grms_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => pc_grms_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => pc_grms_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => pc_grms_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => pc_grms_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => pc_grms_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => pc_grms_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => pc_grms_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => pc_grms_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => pc_grms_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => pc_grms_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => pc_grms_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => pc_grms_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => pc_grms_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => pc_grms_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_007_src_ready,                                                      --              cp.ready
			cp_valid                => cmd_xbar_mux_007_src_valid,                                                      --                .valid
			cp_data                 => cmd_xbar_mux_007_src_data,                                                       --                .data
			cp_startofpacket        => cmd_xbar_mux_007_src_startofpacket,                                              --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_007_src_endofpacket,                                                --                .endofpacket
			cp_channel              => cmd_xbar_mux_007_src_channel,                                                    --                .channel
			rf_sink_ready           => pc_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => pc_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => pc_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => pc_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => pc_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => pc_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => pc_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => pc_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => pc_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => pc_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => pc_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => pc_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => pc_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => pc_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => pc_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => pc_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                            --     (terminated)
			m0_writeresponserequest => open,                                                                            --     (terminated)
			m0_writeresponsevalid   => '0'                                                                              --     (terminated)
		);

	pc_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component p2_grms_qsys_nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 101,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                         --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                  -- clk_reset.reset
			in_data           => pc_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => pc_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => pc_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => pc_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => pc_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => pc_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => pc_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => pc_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => pc_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => pc_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                            -- (terminated)
			csr_read          => '0',                                                                             -- (terminated)
			csr_write         => '0',                                                                             -- (terminated)
			csr_readdata      => open,                                                                            -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                              -- (terminated)
			almost_full_data  => open,                                                                            -- (terminated)
			almost_empty_data => open,                                                                            -- (terminated)
			in_empty          => '0',                                                                             -- (terminated)
			out_empty         => open,                                                                            -- (terminated)
			in_error          => '0',                                                                             -- (terminated)
			out_error         => open,                                                                            -- (terminated)
			in_channel        => '0',                                                                             -- (terminated)
			out_channel       => open                                                                             -- (terminated)
		);

	pd_grms_s1_translator_avalon_universal_slave_0_agent : component p2_grms_qsys_nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 85,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 89,
			PKT_DEST_ID_L             => 86,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 93,
			PKT_PROTECTION_L          => 91,
			PKT_RESPONSE_STATUS_H     => 99,
			PKT_RESPONSE_STATUS_L     => 98,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 14,
			ST_DATA_W                 => 100,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                         --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                  --       clk_reset.reset
			m0_address              => pd_grms_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => pd_grms_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => pd_grms_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => pd_grms_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => pd_grms_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => pd_grms_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => pd_grms_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => pd_grms_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => pd_grms_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => pd_grms_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => pd_grms_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => pd_grms_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => pd_grms_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => pd_grms_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => pd_grms_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => pd_grms_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_008_src_ready,                                                      --              cp.ready
			cp_valid                => cmd_xbar_mux_008_src_valid,                                                      --                .valid
			cp_data                 => cmd_xbar_mux_008_src_data,                                                       --                .data
			cp_startofpacket        => cmd_xbar_mux_008_src_startofpacket,                                              --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_008_src_endofpacket,                                                --                .endofpacket
			cp_channel              => cmd_xbar_mux_008_src_channel,                                                    --                .channel
			rf_sink_ready           => pd_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => pd_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => pd_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => pd_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => pd_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => pd_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => pd_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => pd_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => pd_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => pd_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => pd_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => pd_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => pd_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => pd_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => pd_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => pd_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                            --     (terminated)
			m0_writeresponserequest => open,                                                                            --     (terminated)
			m0_writeresponsevalid   => '0'                                                                              --     (terminated)
		);

	pd_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component p2_grms_qsys_nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 101,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                         --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                  -- clk_reset.reset
			in_data           => pd_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => pd_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => pd_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => pd_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => pd_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => pd_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => pd_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => pd_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => pd_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => pd_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                            -- (terminated)
			csr_read          => '0',                                                                             -- (terminated)
			csr_write         => '0',                                                                             -- (terminated)
			csr_readdata      => open,                                                                            -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                              -- (terminated)
			almost_full_data  => open,                                                                            -- (terminated)
			almost_empty_data => open,                                                                            -- (terminated)
			in_empty          => '0',                                                                             -- (terminated)
			out_empty         => open,                                                                            -- (terminated)
			in_error          => '0',                                                                             -- (terminated)
			out_error         => open,                                                                            -- (terminated)
			in_channel        => '0',                                                                             -- (terminated)
			out_channel       => open                                                                             -- (terminated)
		);

	pe_grms_s1_translator_avalon_universal_slave_0_agent : component p2_grms_qsys_nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 85,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 89,
			PKT_DEST_ID_L             => 86,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 93,
			PKT_PROTECTION_L          => 91,
			PKT_RESPONSE_STATUS_H     => 99,
			PKT_RESPONSE_STATUS_L     => 98,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 14,
			ST_DATA_W                 => 100,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                         --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                  --       clk_reset.reset
			m0_address              => pe_grms_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => pe_grms_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => pe_grms_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => pe_grms_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => pe_grms_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => pe_grms_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => pe_grms_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => pe_grms_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => pe_grms_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => pe_grms_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => pe_grms_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => pe_grms_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => pe_grms_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => pe_grms_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => pe_grms_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => pe_grms_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_009_src_ready,                                                      --              cp.ready
			cp_valid                => cmd_xbar_mux_009_src_valid,                                                      --                .valid
			cp_data                 => cmd_xbar_mux_009_src_data,                                                       --                .data
			cp_startofpacket        => cmd_xbar_mux_009_src_startofpacket,                                              --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_009_src_endofpacket,                                                --                .endofpacket
			cp_channel              => cmd_xbar_mux_009_src_channel,                                                    --                .channel
			rf_sink_ready           => pe_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => pe_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => pe_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => pe_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => pe_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => pe_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => pe_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => pe_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => pe_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => pe_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => pe_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => pe_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => pe_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => pe_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => pe_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => pe_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                            --     (terminated)
			m0_writeresponserequest => open,                                                                            --     (terminated)
			m0_writeresponsevalid   => '0'                                                                              --     (terminated)
		);

	pe_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component p2_grms_qsys_nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 101,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                         --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                  -- clk_reset.reset
			in_data           => pe_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => pe_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => pe_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => pe_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => pe_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => pe_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => pe_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => pe_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => pe_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => pe_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                            -- (terminated)
			csr_read          => '0',                                                                             -- (terminated)
			csr_write         => '0',                                                                             -- (terminated)
			csr_readdata      => open,                                                                            -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                              -- (terminated)
			almost_full_data  => open,                                                                            -- (terminated)
			almost_empty_data => open,                                                                            -- (terminated)
			in_empty          => '0',                                                                             -- (terminated)
			out_empty         => open,                                                                            -- (terminated)
			in_error          => '0',                                                                             -- (terminated)
			out_error         => open,                                                                            -- (terminated)
			in_channel        => '0',                                                                             -- (terminated)
			out_channel       => open                                                                             -- (terminated)
		);

	pf_grms_s1_translator_avalon_universal_slave_0_agent : component p2_grms_qsys_nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 85,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 89,
			PKT_DEST_ID_L             => 86,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 93,
			PKT_PROTECTION_L          => 91,
			PKT_RESPONSE_STATUS_H     => 99,
			PKT_RESPONSE_STATUS_L     => 98,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 14,
			ST_DATA_W                 => 100,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                         --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                  --       clk_reset.reset
			m0_address              => pf_grms_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => pf_grms_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => pf_grms_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => pf_grms_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => pf_grms_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => pf_grms_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => pf_grms_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => pf_grms_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => pf_grms_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => pf_grms_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => pf_grms_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => pf_grms_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => pf_grms_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => pf_grms_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => pf_grms_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => pf_grms_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_010_src_ready,                                                      --              cp.ready
			cp_valid                => cmd_xbar_mux_010_src_valid,                                                      --                .valid
			cp_data                 => cmd_xbar_mux_010_src_data,                                                       --                .data
			cp_startofpacket        => cmd_xbar_mux_010_src_startofpacket,                                              --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_010_src_endofpacket,                                                --                .endofpacket
			cp_channel              => cmd_xbar_mux_010_src_channel,                                                    --                .channel
			rf_sink_ready           => pf_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => pf_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => pf_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => pf_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => pf_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => pf_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => pf_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => pf_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => pf_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => pf_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => pf_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => pf_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => pf_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => pf_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => pf_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => pf_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                            --     (terminated)
			m0_writeresponserequest => open,                                                                            --     (terminated)
			m0_writeresponsevalid   => '0'                                                                              --     (terminated)
		);

	pf_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component p2_grms_qsys_nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 101,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                         --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                  -- clk_reset.reset
			in_data           => pf_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => pf_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => pf_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => pf_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => pf_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => pf_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => pf_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => pf_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => pf_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => pf_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                            -- (terminated)
			csr_read          => '0',                                                                             -- (terminated)
			csr_write         => '0',                                                                             -- (terminated)
			csr_readdata      => open,                                                                            -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                              -- (terminated)
			almost_full_data  => open,                                                                            -- (terminated)
			almost_empty_data => open,                                                                            -- (terminated)
			in_empty          => '0',                                                                             -- (terminated)
			out_empty         => open,                                                                            -- (terminated)
			in_error          => '0',                                                                             -- (terminated)
			out_error         => open,                                                                            -- (terminated)
			in_channel        => '0',                                                                             -- (terminated)
			out_channel       => open                                                                             -- (terminated)
		);

	pg_grms_s1_translator_avalon_universal_slave_0_agent : component p2_grms_qsys_nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 85,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 89,
			PKT_DEST_ID_L             => 86,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 93,
			PKT_PROTECTION_L          => 91,
			PKT_RESPONSE_STATUS_H     => 99,
			PKT_RESPONSE_STATUS_L     => 98,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 14,
			ST_DATA_W                 => 100,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                         --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                  --       clk_reset.reset
			m0_address              => pg_grms_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => pg_grms_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => pg_grms_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => pg_grms_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => pg_grms_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => pg_grms_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => pg_grms_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => pg_grms_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => pg_grms_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => pg_grms_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => pg_grms_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => pg_grms_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => pg_grms_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => pg_grms_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => pg_grms_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => pg_grms_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_011_src_ready,                                                      --              cp.ready
			cp_valid                => cmd_xbar_mux_011_src_valid,                                                      --                .valid
			cp_data                 => cmd_xbar_mux_011_src_data,                                                       --                .data
			cp_startofpacket        => cmd_xbar_mux_011_src_startofpacket,                                              --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_011_src_endofpacket,                                                --                .endofpacket
			cp_channel              => cmd_xbar_mux_011_src_channel,                                                    --                .channel
			rf_sink_ready           => pg_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => pg_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => pg_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => pg_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => pg_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => pg_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => pg_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => pg_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => pg_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => pg_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => pg_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => pg_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => pg_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => pg_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => pg_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => pg_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                            --     (terminated)
			m0_writeresponserequest => open,                                                                            --     (terminated)
			m0_writeresponsevalid   => '0'                                                                              --     (terminated)
		);

	pg_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component p2_grms_qsys_nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 101,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                         --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                  -- clk_reset.reset
			in_data           => pg_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => pg_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => pg_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => pg_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => pg_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => pg_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => pg_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => pg_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => pg_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => pg_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                            -- (terminated)
			csr_read          => '0',                                                                             -- (terminated)
			csr_write         => '0',                                                                             -- (terminated)
			csr_readdata      => open,                                                                            -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                              -- (terminated)
			almost_full_data  => open,                                                                            -- (terminated)
			almost_empty_data => open,                                                                            -- (terminated)
			in_empty          => '0',                                                                             -- (terminated)
			out_empty         => open,                                                                            -- (terminated)
			in_error          => '0',                                                                             -- (terminated)
			out_error         => open,                                                                            -- (terminated)
			in_channel        => '0',                                                                             -- (terminated)
			out_channel       => open                                                                             -- (terminated)
		);

	ph_grms_s1_translator_avalon_universal_slave_0_agent : component p2_grms_qsys_nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 85,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 89,
			PKT_DEST_ID_L             => 86,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 93,
			PKT_PROTECTION_L          => 91,
			PKT_RESPONSE_STATUS_H     => 99,
			PKT_RESPONSE_STATUS_L     => 98,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 14,
			ST_DATA_W                 => 100,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                         --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                  --       clk_reset.reset
			m0_address              => ph_grms_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => ph_grms_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => ph_grms_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => ph_grms_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => ph_grms_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => ph_grms_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => ph_grms_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => ph_grms_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => ph_grms_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => ph_grms_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => ph_grms_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => ph_grms_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => ph_grms_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => ph_grms_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => ph_grms_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => ph_grms_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_012_src_ready,                                                      --              cp.ready
			cp_valid                => cmd_xbar_mux_012_src_valid,                                                      --                .valid
			cp_data                 => cmd_xbar_mux_012_src_data,                                                       --                .data
			cp_startofpacket        => cmd_xbar_mux_012_src_startofpacket,                                              --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_012_src_endofpacket,                                                --                .endofpacket
			cp_channel              => cmd_xbar_mux_012_src_channel,                                                    --                .channel
			rf_sink_ready           => ph_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => ph_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => ph_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => ph_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => ph_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => ph_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => ph_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => ph_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => ph_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => ph_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => ph_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => ph_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => ph_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => ph_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => ph_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => ph_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                            --     (terminated)
			m0_writeresponserequest => open,                                                                            --     (terminated)
			m0_writeresponsevalid   => '0'                                                                              --     (terminated)
		);

	ph_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component p2_grms_qsys_nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 101,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                         --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                  -- clk_reset.reset
			in_data           => ph_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => ph_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => ph_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => ph_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => ph_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => ph_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => ph_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => ph_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => ph_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => ph_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                            -- (terminated)
			csr_read          => '0',                                                                             -- (terminated)
			csr_write         => '0',                                                                             -- (terminated)
			csr_readdata      => open,                                                                            -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                              -- (terminated)
			almost_full_data  => open,                                                                            -- (terminated)
			almost_empty_data => open,                                                                            -- (terminated)
			in_empty          => '0',                                                                             -- (terminated)
			out_empty         => open,                                                                            -- (terminated)
			in_error          => '0',                                                                             -- (terminated)
			out_error         => open,                                                                            -- (terminated)
			in_channel        => '0',                                                                             -- (terminated)
			out_channel       => open                                                                             -- (terminated)
		);

	pi_grms_s1_translator_avalon_universal_slave_0_agent : component p2_grms_qsys_nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 85,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 89,
			PKT_DEST_ID_L             => 86,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 93,
			PKT_PROTECTION_L          => 91,
			PKT_RESPONSE_STATUS_H     => 99,
			PKT_RESPONSE_STATUS_L     => 98,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 14,
			ST_DATA_W                 => 100,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                         --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                  --       clk_reset.reset
			m0_address              => pi_grms_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => pi_grms_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => pi_grms_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => pi_grms_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => pi_grms_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => pi_grms_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => pi_grms_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => pi_grms_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => pi_grms_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => pi_grms_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => pi_grms_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => pi_grms_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => pi_grms_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => pi_grms_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => pi_grms_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => pi_grms_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_013_src_ready,                                                      --              cp.ready
			cp_valid                => cmd_xbar_mux_013_src_valid,                                                      --                .valid
			cp_data                 => cmd_xbar_mux_013_src_data,                                                       --                .data
			cp_startofpacket        => cmd_xbar_mux_013_src_startofpacket,                                              --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_013_src_endofpacket,                                                --                .endofpacket
			cp_channel              => cmd_xbar_mux_013_src_channel,                                                    --                .channel
			rf_sink_ready           => pi_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => pi_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => pi_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => pi_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => pi_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => pi_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => pi_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => pi_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => pi_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => pi_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => pi_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => pi_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => pi_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => pi_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => pi_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => pi_grms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                            --     (terminated)
			m0_writeresponserequest => open,                                                                            --     (terminated)
			m0_writeresponsevalid   => '0'                                                                              --     (terminated)
		);

	pi_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component p2_grms_qsys_nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 101,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                         --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                  -- clk_reset.reset
			in_data           => pi_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => pi_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => pi_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => pi_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => pi_grms_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => pi_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => pi_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => pi_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => pi_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => pi_grms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                            -- (terminated)
			csr_read          => '0',                                                                             -- (terminated)
			csr_write         => '0',                                                                             -- (terminated)
			csr_readdata      => open,                                                                            -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                              -- (terminated)
			almost_full_data  => open,                                                                            -- (terminated)
			almost_empty_data => open,                                                                            -- (terminated)
			in_empty          => '0',                                                                             -- (terminated)
			out_empty         => open,                                                                            -- (terminated)
			in_error          => '0',                                                                             -- (terminated)
			out_error         => open,                                                                            -- (terminated)
			in_channel        => '0',                                                                             -- (terminated)
			out_channel       => open                                                                             -- (terminated)
		);

	addr_router : component p2_grms_qsys_addr_router
		port map (
			sink_ready         => nios2_qsys_grms_instruction_master_translator_avalon_universal_master_0_agent_cp_ready,         --      sink.ready
			sink_valid         => nios2_qsys_grms_instruction_master_translator_avalon_universal_master_0_agent_cp_valid,         --          .valid
			sink_data          => nios2_qsys_grms_instruction_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			sink_startofpacket => nios2_qsys_grms_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			sink_endofpacket   => nios2_qsys_grms_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                                        --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                                 -- clk_reset.reset
			src_ready          => addr_router_src_ready,                                                                          --       src.ready
			src_valid          => addr_router_src_valid,                                                                          --          .valid
			src_data           => addr_router_src_data,                                                                           --          .data
			src_channel        => addr_router_src_channel,                                                                        --          .channel
			src_startofpacket  => addr_router_src_startofpacket,                                                                  --          .startofpacket
			src_endofpacket    => addr_router_src_endofpacket                                                                     --          .endofpacket
		);

	addr_router_001 : component p2_grms_qsys_addr_router
		port map (
			sink_ready         => nios2_qsys_grms_data_master_translator_avalon_universal_master_0_agent_cp_ready,         --      sink.ready
			sink_valid         => nios2_qsys_grms_data_master_translator_avalon_universal_master_0_agent_cp_valid,         --          .valid
			sink_data          => nios2_qsys_grms_data_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			sink_startofpacket => nios2_qsys_grms_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			sink_endofpacket   => nios2_qsys_grms_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                                 --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                          -- clk_reset.reset
			src_ready          => addr_router_001_src_ready,                                                               --       src.ready
			src_valid          => addr_router_001_src_valid,                                                               --          .valid
			src_data           => addr_router_001_src_data,                                                                --          .data
			src_channel        => addr_router_001_src_channel,                                                             --          .channel
			src_startofpacket  => addr_router_001_src_startofpacket,                                                       --          .startofpacket
			src_endofpacket    => addr_router_001_src_endofpacket                                                          --          .endofpacket
		);

	id_router : component p2_grms_qsys_id_router
		port map (
			sink_ready         => nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => nios2_qsys_grms_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                                      --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                               -- clk_reset.reset
			src_ready          => id_router_src_ready,                                                                          --       src.ready
			src_valid          => id_router_src_valid,                                                                          --          .valid
			src_data           => id_router_src_data,                                                                           --          .data
			src_channel        => id_router_src_channel,                                                                        --          .channel
			src_startofpacket  => id_router_src_startofpacket,                                                                  --          .startofpacket
			src_endofpacket    => id_router_src_endofpacket                                                                     --          .endofpacket
		);

	id_router_001 : component p2_grms_qsys_id_router
		port map (
			sink_ready         => jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => jtag_uart_grms_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                                     --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                              -- clk_reset.reset
			src_ready          => id_router_001_src_ready,                                                                     --       src.ready
			src_valid          => id_router_001_src_valid,                                                                     --          .valid
			src_data           => id_router_001_src_data,                                                                      --          .data
			src_channel        => id_router_001_src_channel,                                                                   --          .channel
			src_startofpacket  => id_router_001_src_startofpacket,                                                             --          .startofpacket
			src_endofpacket    => id_router_001_src_endofpacket                                                                --          .endofpacket
		);

	id_router_002 : component p2_grms_qsys_id_router_002
		port map (
			sink_ready         => new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => new_sdram_controller_grms_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                                 --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                          -- clk_reset.reset
			src_ready          => id_router_002_src_ready,                                                                 --       src.ready
			src_valid          => id_router_002_src_valid,                                                                 --          .valid
			src_data           => id_router_002_src_data,                                                                  --          .data
			src_channel        => id_router_002_src_channel,                                                               --          .channel
			src_startofpacket  => id_router_002_src_startofpacket,                                                         --          .startofpacket
			src_endofpacket    => id_router_002_src_endofpacket                                                            --          .endofpacket
		);

	id_router_003 : component p2_grms_qsys_id_router
		port map (
			sink_ready         => timer_grms_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => timer_grms_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => timer_grms_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => timer_grms_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => timer_grms_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                  --       clk.clk
			reset              => rst_controller_reset_out_reset,                                           -- clk_reset.reset
			src_ready          => id_router_003_src_ready,                                                  --       src.ready
			src_valid          => id_router_003_src_valid,                                                  --          .valid
			src_data           => id_router_003_src_data,                                                   --          .data
			src_channel        => id_router_003_src_channel,                                                --          .channel
			src_startofpacket  => id_router_003_src_startofpacket,                                          --          .startofpacket
			src_endofpacket    => id_router_003_src_endofpacket                                             --          .endofpacket
		);

	id_router_004 : component p2_grms_qsys_id_router
		port map (
			sink_ready         => lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => lcd_16207_grms_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                                 --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                          -- clk_reset.reset
			src_ready          => id_router_004_src_ready,                                                                 --       src.ready
			src_valid          => id_router_004_src_valid,                                                                 --          .valid
			src_data           => id_router_004_src_data,                                                                  --          .data
			src_channel        => id_router_004_src_channel,                                                               --          .channel
			src_startofpacket  => id_router_004_src_startofpacket,                                                         --          .startofpacket
			src_endofpacket    => id_router_004_src_endofpacket                                                            --          .endofpacket
		);

	id_router_005 : component p2_grms_qsys_id_router
		port map (
			sink_ready         => pa_grms_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => pa_grms_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => pa_grms_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => pa_grms_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => pa_grms_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                               --       clk.clk
			reset              => rst_controller_reset_out_reset,                                        -- clk_reset.reset
			src_ready          => id_router_005_src_ready,                                               --       src.ready
			src_valid          => id_router_005_src_valid,                                               --          .valid
			src_data           => id_router_005_src_data,                                                --          .data
			src_channel        => id_router_005_src_channel,                                             --          .channel
			src_startofpacket  => id_router_005_src_startofpacket,                                       --          .startofpacket
			src_endofpacket    => id_router_005_src_endofpacket                                          --          .endofpacket
		);

	id_router_006 : component p2_grms_qsys_id_router
		port map (
			sink_ready         => pb_grms_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => pb_grms_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => pb_grms_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => pb_grms_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => pb_grms_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                               --       clk.clk
			reset              => rst_controller_reset_out_reset,                                        -- clk_reset.reset
			src_ready          => id_router_006_src_ready,                                               --       src.ready
			src_valid          => id_router_006_src_valid,                                               --          .valid
			src_data           => id_router_006_src_data,                                                --          .data
			src_channel        => id_router_006_src_channel,                                             --          .channel
			src_startofpacket  => id_router_006_src_startofpacket,                                       --          .startofpacket
			src_endofpacket    => id_router_006_src_endofpacket                                          --          .endofpacket
		);

	id_router_007 : component p2_grms_qsys_id_router
		port map (
			sink_ready         => pc_grms_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => pc_grms_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => pc_grms_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => pc_grms_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => pc_grms_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                               --       clk.clk
			reset              => rst_controller_reset_out_reset,                                        -- clk_reset.reset
			src_ready          => id_router_007_src_ready,                                               --       src.ready
			src_valid          => id_router_007_src_valid,                                               --          .valid
			src_data           => id_router_007_src_data,                                                --          .data
			src_channel        => id_router_007_src_channel,                                             --          .channel
			src_startofpacket  => id_router_007_src_startofpacket,                                       --          .startofpacket
			src_endofpacket    => id_router_007_src_endofpacket                                          --          .endofpacket
		);

	id_router_008 : component p2_grms_qsys_id_router
		port map (
			sink_ready         => pd_grms_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => pd_grms_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => pd_grms_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => pd_grms_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => pd_grms_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                               --       clk.clk
			reset              => rst_controller_reset_out_reset,                                        -- clk_reset.reset
			src_ready          => id_router_008_src_ready,                                               --       src.ready
			src_valid          => id_router_008_src_valid,                                               --          .valid
			src_data           => id_router_008_src_data,                                                --          .data
			src_channel        => id_router_008_src_channel,                                             --          .channel
			src_startofpacket  => id_router_008_src_startofpacket,                                       --          .startofpacket
			src_endofpacket    => id_router_008_src_endofpacket                                          --          .endofpacket
		);

	id_router_009 : component p2_grms_qsys_id_router
		port map (
			sink_ready         => pe_grms_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => pe_grms_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => pe_grms_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => pe_grms_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => pe_grms_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                               --       clk.clk
			reset              => rst_controller_reset_out_reset,                                        -- clk_reset.reset
			src_ready          => id_router_009_src_ready,                                               --       src.ready
			src_valid          => id_router_009_src_valid,                                               --          .valid
			src_data           => id_router_009_src_data,                                                --          .data
			src_channel        => id_router_009_src_channel,                                             --          .channel
			src_startofpacket  => id_router_009_src_startofpacket,                                       --          .startofpacket
			src_endofpacket    => id_router_009_src_endofpacket                                          --          .endofpacket
		);

	id_router_010 : component p2_grms_qsys_id_router
		port map (
			sink_ready         => pf_grms_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => pf_grms_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => pf_grms_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => pf_grms_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => pf_grms_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                               --       clk.clk
			reset              => rst_controller_reset_out_reset,                                        -- clk_reset.reset
			src_ready          => id_router_010_src_ready,                                               --       src.ready
			src_valid          => id_router_010_src_valid,                                               --          .valid
			src_data           => id_router_010_src_data,                                                --          .data
			src_channel        => id_router_010_src_channel,                                             --          .channel
			src_startofpacket  => id_router_010_src_startofpacket,                                       --          .startofpacket
			src_endofpacket    => id_router_010_src_endofpacket                                          --          .endofpacket
		);

	id_router_011 : component p2_grms_qsys_id_router
		port map (
			sink_ready         => pg_grms_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => pg_grms_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => pg_grms_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => pg_grms_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => pg_grms_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                               --       clk.clk
			reset              => rst_controller_reset_out_reset,                                        -- clk_reset.reset
			src_ready          => id_router_011_src_ready,                                               --       src.ready
			src_valid          => id_router_011_src_valid,                                               --          .valid
			src_data           => id_router_011_src_data,                                                --          .data
			src_channel        => id_router_011_src_channel,                                             --          .channel
			src_startofpacket  => id_router_011_src_startofpacket,                                       --          .startofpacket
			src_endofpacket    => id_router_011_src_endofpacket                                          --          .endofpacket
		);

	id_router_012 : component p2_grms_qsys_id_router
		port map (
			sink_ready         => ph_grms_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => ph_grms_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => ph_grms_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => ph_grms_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => ph_grms_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                               --       clk.clk
			reset              => rst_controller_reset_out_reset,                                        -- clk_reset.reset
			src_ready          => id_router_012_src_ready,                                               --       src.ready
			src_valid          => id_router_012_src_valid,                                               --          .valid
			src_data           => id_router_012_src_data,                                                --          .data
			src_channel        => id_router_012_src_channel,                                             --          .channel
			src_startofpacket  => id_router_012_src_startofpacket,                                       --          .startofpacket
			src_endofpacket    => id_router_012_src_endofpacket                                          --          .endofpacket
		);

	id_router_013 : component p2_grms_qsys_id_router
		port map (
			sink_ready         => pi_grms_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => pi_grms_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => pi_grms_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => pi_grms_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => pi_grms_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                               --       clk.clk
			reset              => rst_controller_reset_out_reset,                                        -- clk_reset.reset
			src_ready          => id_router_013_src_ready,                                               --       src.ready
			src_valid          => id_router_013_src_valid,                                               --          .valid
			src_data           => id_router_013_src_data,                                                --          .data
			src_channel        => id_router_013_src_channel,                                             --          .channel
			src_startofpacket  => id_router_013_src_startofpacket,                                       --          .startofpacket
			src_endofpacket    => id_router_013_src_endofpacket                                          --          .endofpacket
		);

	burst_adapter : component altera_merlin_burst_adapter
		generic map (
			PKT_ADDR_H                => 42,
			PKT_ADDR_L                => 18,
			PKT_BEGIN_BURST           => 62,
			PKT_BYTE_CNT_H            => 51,
			PKT_BYTE_CNT_L            => 49,
			PKT_BYTEEN_H              => 17,
			PKT_BYTEEN_L              => 16,
			PKT_BURST_SIZE_H          => 57,
			PKT_BURST_SIZE_L          => 55,
			PKT_BURST_TYPE_H          => 59,
			PKT_BURST_TYPE_L          => 58,
			PKT_BURSTWRAP_H           => 54,
			PKT_BURSTWRAP_L           => 52,
			PKT_TRANS_COMPRESSED_READ => 43,
			PKT_TRANS_WRITE           => 45,
			PKT_TRANS_READ            => 46,
			OUT_NARROW_SIZE           => 0,
			IN_NARROW_SIZE            => 0,
			OUT_FIXED                 => 0,
			OUT_COMPLETE_WRAP         => 0,
			ST_DATA_W                 => 82,
			ST_CHANNEL_W              => 14,
			OUT_BYTE_CNT_H            => 50,
			OUT_BURSTWRAP_H           => 54,
			COMPRESSED_READ_SUPPORT   => 0,
			BYTEENABLE_SYNTHESIS      => 1,
			PIPE_INPUTS               => 0,
			NO_WRAP_SUPPORT           => 0,
			BURSTWRAP_CONST_MASK      => 3,
			BURSTWRAP_CONST_VALUE     => 3
		)
		port map (
			clk                   => clk_clk,                             --       cr0.clk
			reset                 => rst_controller_reset_out_reset,      -- cr0_reset.reset
			sink0_valid           => width_adapter_src_valid,             --     sink0.valid
			sink0_data            => width_adapter_src_data,              --          .data
			sink0_channel         => width_adapter_src_channel,           --          .channel
			sink0_startofpacket   => width_adapter_src_startofpacket,     --          .startofpacket
			sink0_endofpacket     => width_adapter_src_endofpacket,       --          .endofpacket
			sink0_ready           => width_adapter_src_ready,             --          .ready
			source0_valid         => burst_adapter_source0_valid,         --   source0.valid
			source0_data          => burst_adapter_source0_data,          --          .data
			source0_channel       => burst_adapter_source0_channel,       --          .channel
			source0_startofpacket => burst_adapter_source0_startofpacket, --          .startofpacket
			source0_endofpacket   => burst_adapter_source0_endofpacket,   --          .endofpacket
			source0_ready         => burst_adapter_source0_ready          --          .ready
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS        => 1,
			OUTPUT_RESET_SYNC_EDGES => "deassert",
			SYNC_DEPTH              => 2,
			RESET_REQUEST_PRESENT   => 0
		)
		port map (
			reset_in0  => reset_reset_n_ports_inv,        -- reset_in0.reset
			clk        => clk_clk,                        --       clk.clk
			reset_out  => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req  => open,                           -- (terminated)
			reset_in1  => '0',                            -- (terminated)
			reset_in2  => '0',                            -- (terminated)
			reset_in3  => '0',                            -- (terminated)
			reset_in4  => '0',                            -- (terminated)
			reset_in5  => '0',                            -- (terminated)
			reset_in6  => '0',                            -- (terminated)
			reset_in7  => '0',                            -- (terminated)
			reset_in8  => '0',                            -- (terminated)
			reset_in9  => '0',                            -- (terminated)
			reset_in10 => '0',                            -- (terminated)
			reset_in11 => '0',                            -- (terminated)
			reset_in12 => '0',                            -- (terminated)
			reset_in13 => '0',                            -- (terminated)
			reset_in14 => '0',                            -- (terminated)
			reset_in15 => '0'                             -- (terminated)
		);

	cmd_xbar_demux : component p2_grms_qsys_cmd_xbar_demux
		port map (
			clk                 => clk_clk,                            --       clk.clk
			reset               => rst_controller_reset_out_reset,     -- clk_reset.reset
			sink_ready          => addr_router_src_ready,              --      sink.ready
			sink_channel        => addr_router_src_channel,            --          .channel
			sink_data           => addr_router_src_data,               --          .data
			sink_startofpacket  => addr_router_src_startofpacket,      --          .startofpacket
			sink_endofpacket    => addr_router_src_endofpacket,        --          .endofpacket
			sink_valid(0)       => addr_router_src_valid,              --          .valid
			src0_ready          => cmd_xbar_demux_src0_ready,          --      src0.ready
			src0_valid          => cmd_xbar_demux_src0_valid,          --          .valid
			src0_data           => cmd_xbar_demux_src0_data,           --          .data
			src0_channel        => cmd_xbar_demux_src0_channel,        --          .channel
			src0_startofpacket  => cmd_xbar_demux_src0_startofpacket,  --          .startofpacket
			src0_endofpacket    => cmd_xbar_demux_src0_endofpacket,    --          .endofpacket
			src1_ready          => cmd_xbar_demux_src1_ready,          --      src1.ready
			src1_valid          => cmd_xbar_demux_src1_valid,          --          .valid
			src1_data           => cmd_xbar_demux_src1_data,           --          .data
			src1_channel        => cmd_xbar_demux_src1_channel,        --          .channel
			src1_startofpacket  => cmd_xbar_demux_src1_startofpacket,  --          .startofpacket
			src1_endofpacket    => cmd_xbar_demux_src1_endofpacket,    --          .endofpacket
			src2_ready          => cmd_xbar_demux_src2_ready,          --      src2.ready
			src2_valid          => cmd_xbar_demux_src2_valid,          --          .valid
			src2_data           => cmd_xbar_demux_src2_data,           --          .data
			src2_channel        => cmd_xbar_demux_src2_channel,        --          .channel
			src2_startofpacket  => cmd_xbar_demux_src2_startofpacket,  --          .startofpacket
			src2_endofpacket    => cmd_xbar_demux_src2_endofpacket,    --          .endofpacket
			src3_ready          => cmd_xbar_demux_src3_ready,          --      src3.ready
			src3_valid          => cmd_xbar_demux_src3_valid,          --          .valid
			src3_data           => cmd_xbar_demux_src3_data,           --          .data
			src3_channel        => cmd_xbar_demux_src3_channel,        --          .channel
			src3_startofpacket  => cmd_xbar_demux_src3_startofpacket,  --          .startofpacket
			src3_endofpacket    => cmd_xbar_demux_src3_endofpacket,    --          .endofpacket
			src4_ready          => cmd_xbar_demux_src4_ready,          --      src4.ready
			src4_valid          => cmd_xbar_demux_src4_valid,          --          .valid
			src4_data           => cmd_xbar_demux_src4_data,           --          .data
			src4_channel        => cmd_xbar_demux_src4_channel,        --          .channel
			src4_startofpacket  => cmd_xbar_demux_src4_startofpacket,  --          .startofpacket
			src4_endofpacket    => cmd_xbar_demux_src4_endofpacket,    --          .endofpacket
			src5_ready          => cmd_xbar_demux_src5_ready,          --      src5.ready
			src5_valid          => cmd_xbar_demux_src5_valid,          --          .valid
			src5_data           => cmd_xbar_demux_src5_data,           --          .data
			src5_channel        => cmd_xbar_demux_src5_channel,        --          .channel
			src5_startofpacket  => cmd_xbar_demux_src5_startofpacket,  --          .startofpacket
			src5_endofpacket    => cmd_xbar_demux_src5_endofpacket,    --          .endofpacket
			src6_ready          => cmd_xbar_demux_src6_ready,          --      src6.ready
			src6_valid          => cmd_xbar_demux_src6_valid,          --          .valid
			src6_data           => cmd_xbar_demux_src6_data,           --          .data
			src6_channel        => cmd_xbar_demux_src6_channel,        --          .channel
			src6_startofpacket  => cmd_xbar_demux_src6_startofpacket,  --          .startofpacket
			src6_endofpacket    => cmd_xbar_demux_src6_endofpacket,    --          .endofpacket
			src7_ready          => cmd_xbar_demux_src7_ready,          --      src7.ready
			src7_valid          => cmd_xbar_demux_src7_valid,          --          .valid
			src7_data           => cmd_xbar_demux_src7_data,           --          .data
			src7_channel        => cmd_xbar_demux_src7_channel,        --          .channel
			src7_startofpacket  => cmd_xbar_demux_src7_startofpacket,  --          .startofpacket
			src7_endofpacket    => cmd_xbar_demux_src7_endofpacket,    --          .endofpacket
			src8_ready          => cmd_xbar_demux_src8_ready,          --      src8.ready
			src8_valid          => cmd_xbar_demux_src8_valid,          --          .valid
			src8_data           => cmd_xbar_demux_src8_data,           --          .data
			src8_channel        => cmd_xbar_demux_src8_channel,        --          .channel
			src8_startofpacket  => cmd_xbar_demux_src8_startofpacket,  --          .startofpacket
			src8_endofpacket    => cmd_xbar_demux_src8_endofpacket,    --          .endofpacket
			src9_ready          => cmd_xbar_demux_src9_ready,          --      src9.ready
			src9_valid          => cmd_xbar_demux_src9_valid,          --          .valid
			src9_data           => cmd_xbar_demux_src9_data,           --          .data
			src9_channel        => cmd_xbar_demux_src9_channel,        --          .channel
			src9_startofpacket  => cmd_xbar_demux_src9_startofpacket,  --          .startofpacket
			src9_endofpacket    => cmd_xbar_demux_src9_endofpacket,    --          .endofpacket
			src10_ready         => cmd_xbar_demux_src10_ready,         --     src10.ready
			src10_valid         => cmd_xbar_demux_src10_valid,         --          .valid
			src10_data          => cmd_xbar_demux_src10_data,          --          .data
			src10_channel       => cmd_xbar_demux_src10_channel,       --          .channel
			src10_startofpacket => cmd_xbar_demux_src10_startofpacket, --          .startofpacket
			src10_endofpacket   => cmd_xbar_demux_src10_endofpacket,   --          .endofpacket
			src11_ready         => cmd_xbar_demux_src11_ready,         --     src11.ready
			src11_valid         => cmd_xbar_demux_src11_valid,         --          .valid
			src11_data          => cmd_xbar_demux_src11_data,          --          .data
			src11_channel       => cmd_xbar_demux_src11_channel,       --          .channel
			src11_startofpacket => cmd_xbar_demux_src11_startofpacket, --          .startofpacket
			src11_endofpacket   => cmd_xbar_demux_src11_endofpacket,   --          .endofpacket
			src12_ready         => cmd_xbar_demux_src12_ready,         --     src12.ready
			src12_valid         => cmd_xbar_demux_src12_valid,         --          .valid
			src12_data          => cmd_xbar_demux_src12_data,          --          .data
			src12_channel       => cmd_xbar_demux_src12_channel,       --          .channel
			src12_startofpacket => cmd_xbar_demux_src12_startofpacket, --          .startofpacket
			src12_endofpacket   => cmd_xbar_demux_src12_endofpacket,   --          .endofpacket
			src13_ready         => cmd_xbar_demux_src13_ready,         --     src13.ready
			src13_valid         => cmd_xbar_demux_src13_valid,         --          .valid
			src13_data          => cmd_xbar_demux_src13_data,          --          .data
			src13_channel       => cmd_xbar_demux_src13_channel,       --          .channel
			src13_startofpacket => cmd_xbar_demux_src13_startofpacket, --          .startofpacket
			src13_endofpacket   => cmd_xbar_demux_src13_endofpacket    --          .endofpacket
		);

	cmd_xbar_demux_001 : component p2_grms_qsys_cmd_xbar_demux
		port map (
			clk                 => clk_clk,                                --       clk.clk
			reset               => rst_controller_reset_out_reset,         -- clk_reset.reset
			sink_ready          => addr_router_001_src_ready,              --      sink.ready
			sink_channel        => addr_router_001_src_channel,            --          .channel
			sink_data           => addr_router_001_src_data,               --          .data
			sink_startofpacket  => addr_router_001_src_startofpacket,      --          .startofpacket
			sink_endofpacket    => addr_router_001_src_endofpacket,        --          .endofpacket
			sink_valid(0)       => addr_router_001_src_valid,              --          .valid
			src0_ready          => cmd_xbar_demux_001_src0_ready,          --      src0.ready
			src0_valid          => cmd_xbar_demux_001_src0_valid,          --          .valid
			src0_data           => cmd_xbar_demux_001_src0_data,           --          .data
			src0_channel        => cmd_xbar_demux_001_src0_channel,        --          .channel
			src0_startofpacket  => cmd_xbar_demux_001_src0_startofpacket,  --          .startofpacket
			src0_endofpacket    => cmd_xbar_demux_001_src0_endofpacket,    --          .endofpacket
			src1_ready          => cmd_xbar_demux_001_src1_ready,          --      src1.ready
			src1_valid          => cmd_xbar_demux_001_src1_valid,          --          .valid
			src1_data           => cmd_xbar_demux_001_src1_data,           --          .data
			src1_channel        => cmd_xbar_demux_001_src1_channel,        --          .channel
			src1_startofpacket  => cmd_xbar_demux_001_src1_startofpacket,  --          .startofpacket
			src1_endofpacket    => cmd_xbar_demux_001_src1_endofpacket,    --          .endofpacket
			src2_ready          => cmd_xbar_demux_001_src2_ready,          --      src2.ready
			src2_valid          => cmd_xbar_demux_001_src2_valid,          --          .valid
			src2_data           => cmd_xbar_demux_001_src2_data,           --          .data
			src2_channel        => cmd_xbar_demux_001_src2_channel,        --          .channel
			src2_startofpacket  => cmd_xbar_demux_001_src2_startofpacket,  --          .startofpacket
			src2_endofpacket    => cmd_xbar_demux_001_src2_endofpacket,    --          .endofpacket
			src3_ready          => cmd_xbar_demux_001_src3_ready,          --      src3.ready
			src3_valid          => cmd_xbar_demux_001_src3_valid,          --          .valid
			src3_data           => cmd_xbar_demux_001_src3_data,           --          .data
			src3_channel        => cmd_xbar_demux_001_src3_channel,        --          .channel
			src3_startofpacket  => cmd_xbar_demux_001_src3_startofpacket,  --          .startofpacket
			src3_endofpacket    => cmd_xbar_demux_001_src3_endofpacket,    --          .endofpacket
			src4_ready          => cmd_xbar_demux_001_src4_ready,          --      src4.ready
			src4_valid          => cmd_xbar_demux_001_src4_valid,          --          .valid
			src4_data           => cmd_xbar_demux_001_src4_data,           --          .data
			src4_channel        => cmd_xbar_demux_001_src4_channel,        --          .channel
			src4_startofpacket  => cmd_xbar_demux_001_src4_startofpacket,  --          .startofpacket
			src4_endofpacket    => cmd_xbar_demux_001_src4_endofpacket,    --          .endofpacket
			src5_ready          => cmd_xbar_demux_001_src5_ready,          --      src5.ready
			src5_valid          => cmd_xbar_demux_001_src5_valid,          --          .valid
			src5_data           => cmd_xbar_demux_001_src5_data,           --          .data
			src5_channel        => cmd_xbar_demux_001_src5_channel,        --          .channel
			src5_startofpacket  => cmd_xbar_demux_001_src5_startofpacket,  --          .startofpacket
			src5_endofpacket    => cmd_xbar_demux_001_src5_endofpacket,    --          .endofpacket
			src6_ready          => cmd_xbar_demux_001_src6_ready,          --      src6.ready
			src6_valid          => cmd_xbar_demux_001_src6_valid,          --          .valid
			src6_data           => cmd_xbar_demux_001_src6_data,           --          .data
			src6_channel        => cmd_xbar_demux_001_src6_channel,        --          .channel
			src6_startofpacket  => cmd_xbar_demux_001_src6_startofpacket,  --          .startofpacket
			src6_endofpacket    => cmd_xbar_demux_001_src6_endofpacket,    --          .endofpacket
			src7_ready          => cmd_xbar_demux_001_src7_ready,          --      src7.ready
			src7_valid          => cmd_xbar_demux_001_src7_valid,          --          .valid
			src7_data           => cmd_xbar_demux_001_src7_data,           --          .data
			src7_channel        => cmd_xbar_demux_001_src7_channel,        --          .channel
			src7_startofpacket  => cmd_xbar_demux_001_src7_startofpacket,  --          .startofpacket
			src7_endofpacket    => cmd_xbar_demux_001_src7_endofpacket,    --          .endofpacket
			src8_ready          => cmd_xbar_demux_001_src8_ready,          --      src8.ready
			src8_valid          => cmd_xbar_demux_001_src8_valid,          --          .valid
			src8_data           => cmd_xbar_demux_001_src8_data,           --          .data
			src8_channel        => cmd_xbar_demux_001_src8_channel,        --          .channel
			src8_startofpacket  => cmd_xbar_demux_001_src8_startofpacket,  --          .startofpacket
			src8_endofpacket    => cmd_xbar_demux_001_src8_endofpacket,    --          .endofpacket
			src9_ready          => cmd_xbar_demux_001_src9_ready,          --      src9.ready
			src9_valid          => cmd_xbar_demux_001_src9_valid,          --          .valid
			src9_data           => cmd_xbar_demux_001_src9_data,           --          .data
			src9_channel        => cmd_xbar_demux_001_src9_channel,        --          .channel
			src9_startofpacket  => cmd_xbar_demux_001_src9_startofpacket,  --          .startofpacket
			src9_endofpacket    => cmd_xbar_demux_001_src9_endofpacket,    --          .endofpacket
			src10_ready         => cmd_xbar_demux_001_src10_ready,         --     src10.ready
			src10_valid         => cmd_xbar_demux_001_src10_valid,         --          .valid
			src10_data          => cmd_xbar_demux_001_src10_data,          --          .data
			src10_channel       => cmd_xbar_demux_001_src10_channel,       --          .channel
			src10_startofpacket => cmd_xbar_demux_001_src10_startofpacket, --          .startofpacket
			src10_endofpacket   => cmd_xbar_demux_001_src10_endofpacket,   --          .endofpacket
			src11_ready         => cmd_xbar_demux_001_src11_ready,         --     src11.ready
			src11_valid         => cmd_xbar_demux_001_src11_valid,         --          .valid
			src11_data          => cmd_xbar_demux_001_src11_data,          --          .data
			src11_channel       => cmd_xbar_demux_001_src11_channel,       --          .channel
			src11_startofpacket => cmd_xbar_demux_001_src11_startofpacket, --          .startofpacket
			src11_endofpacket   => cmd_xbar_demux_001_src11_endofpacket,   --          .endofpacket
			src12_ready         => cmd_xbar_demux_001_src12_ready,         --     src12.ready
			src12_valid         => cmd_xbar_demux_001_src12_valid,         --          .valid
			src12_data          => cmd_xbar_demux_001_src12_data,          --          .data
			src12_channel       => cmd_xbar_demux_001_src12_channel,       --          .channel
			src12_startofpacket => cmd_xbar_demux_001_src12_startofpacket, --          .startofpacket
			src12_endofpacket   => cmd_xbar_demux_001_src12_endofpacket,   --          .endofpacket
			src13_ready         => cmd_xbar_demux_001_src13_ready,         --     src13.ready
			src13_valid         => cmd_xbar_demux_001_src13_valid,         --          .valid
			src13_data          => cmd_xbar_demux_001_src13_data,          --          .data
			src13_channel       => cmd_xbar_demux_001_src13_channel,       --          .channel
			src13_startofpacket => cmd_xbar_demux_001_src13_startofpacket, --          .startofpacket
			src13_endofpacket   => cmd_xbar_demux_001_src13_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux : component p2_grms_qsys_cmd_xbar_mux
		port map (
			clk                 => clk_clk,                               --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => cmd_xbar_mux_src_ready,                --       src.ready
			src_valid           => cmd_xbar_mux_src_valid,                --          .valid
			src_data            => cmd_xbar_mux_src_data,                 --          .data
			src_channel         => cmd_xbar_mux_src_channel,              --          .channel
			src_startofpacket   => cmd_xbar_mux_src_startofpacket,        --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_src_endofpacket,          --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src0_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src0_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src0_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src0_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src0_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src0_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src0_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src0_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src0_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src0_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src0_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src0_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_001 : component p2_grms_qsys_cmd_xbar_mux
		port map (
			clk                 => clk_clk,                               --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => cmd_xbar_mux_001_src_ready,            --       src.ready
			src_valid           => cmd_xbar_mux_001_src_valid,            --          .valid
			src_data            => cmd_xbar_mux_001_src_data,             --          .data
			src_channel         => cmd_xbar_mux_001_src_channel,          --          .channel
			src_startofpacket   => cmd_xbar_mux_001_src_startofpacket,    --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_001_src_endofpacket,      --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src1_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src1_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src1_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src1_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src1_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src1_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src1_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src1_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src1_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src1_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src1_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src1_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_002 : component p2_grms_qsys_cmd_xbar_mux
		port map (
			clk                 => clk_clk,                               --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => cmd_xbar_mux_002_src_ready,            --       src.ready
			src_valid           => cmd_xbar_mux_002_src_valid,            --          .valid
			src_data            => cmd_xbar_mux_002_src_data,             --          .data
			src_channel         => cmd_xbar_mux_002_src_channel,          --          .channel
			src_startofpacket   => cmd_xbar_mux_002_src_startofpacket,    --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_002_src_endofpacket,      --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src2_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src2_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src2_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src2_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src2_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src2_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src2_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src2_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src2_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src2_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src2_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src2_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_003 : component p2_grms_qsys_cmd_xbar_mux
		port map (
			clk                 => clk_clk,                               --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => cmd_xbar_mux_003_src_ready,            --       src.ready
			src_valid           => cmd_xbar_mux_003_src_valid,            --          .valid
			src_data            => cmd_xbar_mux_003_src_data,             --          .data
			src_channel         => cmd_xbar_mux_003_src_channel,          --          .channel
			src_startofpacket   => cmd_xbar_mux_003_src_startofpacket,    --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_003_src_endofpacket,      --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src3_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src3_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src3_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src3_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src3_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src3_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src3_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src3_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src3_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src3_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src3_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src3_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_004 : component p2_grms_qsys_cmd_xbar_mux
		port map (
			clk                 => clk_clk,                               --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => cmd_xbar_mux_004_src_ready,            --       src.ready
			src_valid           => cmd_xbar_mux_004_src_valid,            --          .valid
			src_data            => cmd_xbar_mux_004_src_data,             --          .data
			src_channel         => cmd_xbar_mux_004_src_channel,          --          .channel
			src_startofpacket   => cmd_xbar_mux_004_src_startofpacket,    --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_004_src_endofpacket,      --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src4_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src4_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src4_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src4_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src4_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src4_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src4_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src4_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src4_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src4_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src4_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src4_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_005 : component p2_grms_qsys_cmd_xbar_mux
		port map (
			clk                 => clk_clk,                               --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => cmd_xbar_mux_005_src_ready,            --       src.ready
			src_valid           => cmd_xbar_mux_005_src_valid,            --          .valid
			src_data            => cmd_xbar_mux_005_src_data,             --          .data
			src_channel         => cmd_xbar_mux_005_src_channel,          --          .channel
			src_startofpacket   => cmd_xbar_mux_005_src_startofpacket,    --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_005_src_endofpacket,      --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src5_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src5_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src5_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src5_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src5_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src5_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src5_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src5_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src5_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src5_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src5_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src5_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_006 : component p2_grms_qsys_cmd_xbar_mux
		port map (
			clk                 => clk_clk,                               --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => cmd_xbar_mux_006_src_ready,            --       src.ready
			src_valid           => cmd_xbar_mux_006_src_valid,            --          .valid
			src_data            => cmd_xbar_mux_006_src_data,             --          .data
			src_channel         => cmd_xbar_mux_006_src_channel,          --          .channel
			src_startofpacket   => cmd_xbar_mux_006_src_startofpacket,    --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_006_src_endofpacket,      --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src6_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src6_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src6_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src6_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src6_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src6_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src6_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src6_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src6_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src6_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src6_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src6_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_007 : component p2_grms_qsys_cmd_xbar_mux
		port map (
			clk                 => clk_clk,                               --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => cmd_xbar_mux_007_src_ready,            --       src.ready
			src_valid           => cmd_xbar_mux_007_src_valid,            --          .valid
			src_data            => cmd_xbar_mux_007_src_data,             --          .data
			src_channel         => cmd_xbar_mux_007_src_channel,          --          .channel
			src_startofpacket   => cmd_xbar_mux_007_src_startofpacket,    --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_007_src_endofpacket,      --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src7_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src7_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src7_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src7_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src7_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src7_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src7_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src7_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src7_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src7_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src7_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src7_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_008 : component p2_grms_qsys_cmd_xbar_mux
		port map (
			clk                 => clk_clk,                               --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => cmd_xbar_mux_008_src_ready,            --       src.ready
			src_valid           => cmd_xbar_mux_008_src_valid,            --          .valid
			src_data            => cmd_xbar_mux_008_src_data,             --          .data
			src_channel         => cmd_xbar_mux_008_src_channel,          --          .channel
			src_startofpacket   => cmd_xbar_mux_008_src_startofpacket,    --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_008_src_endofpacket,      --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src8_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src8_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src8_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src8_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src8_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src8_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src8_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src8_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src8_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src8_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src8_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src8_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_009 : component p2_grms_qsys_cmd_xbar_mux
		port map (
			clk                 => clk_clk,                               --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => cmd_xbar_mux_009_src_ready,            --       src.ready
			src_valid           => cmd_xbar_mux_009_src_valid,            --          .valid
			src_data            => cmd_xbar_mux_009_src_data,             --          .data
			src_channel         => cmd_xbar_mux_009_src_channel,          --          .channel
			src_startofpacket   => cmd_xbar_mux_009_src_startofpacket,    --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_009_src_endofpacket,      --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src9_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src9_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src9_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src9_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src9_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src9_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src9_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src9_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src9_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src9_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src9_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src9_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_010 : component p2_grms_qsys_cmd_xbar_mux
		port map (
			clk                 => clk_clk,                                --       clk.clk
			reset               => rst_controller_reset_out_reset,         -- clk_reset.reset
			src_ready           => cmd_xbar_mux_010_src_ready,             --       src.ready
			src_valid           => cmd_xbar_mux_010_src_valid,             --          .valid
			src_data            => cmd_xbar_mux_010_src_data,              --          .data
			src_channel         => cmd_xbar_mux_010_src_channel,           --          .channel
			src_startofpacket   => cmd_xbar_mux_010_src_startofpacket,     --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_010_src_endofpacket,       --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src10_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src10_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src10_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src10_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src10_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src10_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src10_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src10_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src10_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src10_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src10_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src10_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_011 : component p2_grms_qsys_cmd_xbar_mux
		port map (
			clk                 => clk_clk,                                --       clk.clk
			reset               => rst_controller_reset_out_reset,         -- clk_reset.reset
			src_ready           => cmd_xbar_mux_011_src_ready,             --       src.ready
			src_valid           => cmd_xbar_mux_011_src_valid,             --          .valid
			src_data            => cmd_xbar_mux_011_src_data,              --          .data
			src_channel         => cmd_xbar_mux_011_src_channel,           --          .channel
			src_startofpacket   => cmd_xbar_mux_011_src_startofpacket,     --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_011_src_endofpacket,       --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src11_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src11_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src11_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src11_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src11_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src11_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src11_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src11_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src11_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src11_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src11_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src11_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_012 : component p2_grms_qsys_cmd_xbar_mux
		port map (
			clk                 => clk_clk,                                --       clk.clk
			reset               => rst_controller_reset_out_reset,         -- clk_reset.reset
			src_ready           => cmd_xbar_mux_012_src_ready,             --       src.ready
			src_valid           => cmd_xbar_mux_012_src_valid,             --          .valid
			src_data            => cmd_xbar_mux_012_src_data,              --          .data
			src_channel         => cmd_xbar_mux_012_src_channel,           --          .channel
			src_startofpacket   => cmd_xbar_mux_012_src_startofpacket,     --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_012_src_endofpacket,       --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src12_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src12_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src12_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src12_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src12_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src12_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src12_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src12_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src12_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src12_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src12_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src12_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_013 : component p2_grms_qsys_cmd_xbar_mux
		port map (
			clk                 => clk_clk,                                --       clk.clk
			reset               => rst_controller_reset_out_reset,         -- clk_reset.reset
			src_ready           => cmd_xbar_mux_013_src_ready,             --       src.ready
			src_valid           => cmd_xbar_mux_013_src_valid,             --          .valid
			src_data            => cmd_xbar_mux_013_src_data,              --          .data
			src_channel         => cmd_xbar_mux_013_src_channel,           --          .channel
			src_startofpacket   => cmd_xbar_mux_013_src_startofpacket,     --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_013_src_endofpacket,       --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src13_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src13_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src13_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src13_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src13_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src13_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src13_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src13_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src13_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src13_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src13_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src13_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux : component p2_grms_qsys_rsp_xbar_demux
		port map (
			clk                => clk_clk,                           --       clk.clk
			reset              => rst_controller_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_src_ready,               --      sink.ready
			sink_channel       => id_router_src_channel,             --          .channel
			sink_data          => id_router_src_data,                --          .data
			sink_startofpacket => id_router_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_001 : component p2_grms_qsys_rsp_xbar_demux
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_001_src_ready,               --      sink.ready
			sink_channel       => id_router_001_src_channel,             --          .channel
			sink_data          => id_router_001_src_data,                --          .data
			sink_startofpacket => id_router_001_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_001_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_001_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_001_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_001_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_001_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_001_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_001_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_001_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_001_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_001_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_001_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_001_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_001_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_001_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_002 : component p2_grms_qsys_rsp_xbar_demux
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => width_adapter_001_src_ready,           --      sink.ready
			sink_channel       => width_adapter_001_src_channel,         --          .channel
			sink_data          => width_adapter_001_src_data,            --          .data
			sink_startofpacket => width_adapter_001_src_startofpacket,   --          .startofpacket
			sink_endofpacket   => width_adapter_001_src_endofpacket,     --          .endofpacket
			sink_valid(0)      => width_adapter_001_src_valid,           --          .valid
			src0_ready         => rsp_xbar_demux_002_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_002_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_002_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_002_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_002_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_002_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_002_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_002_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_002_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_002_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_002_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_002_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_003 : component p2_grms_qsys_rsp_xbar_demux
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_003_src_ready,               --      sink.ready
			sink_channel       => id_router_003_src_channel,             --          .channel
			sink_data          => id_router_003_src_data,                --          .data
			sink_startofpacket => id_router_003_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_003_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_003_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_003_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_003_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_003_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_003_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_003_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_003_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_003_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_003_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_003_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_003_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_003_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_003_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_004 : component p2_grms_qsys_rsp_xbar_demux
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_004_src_ready,               --      sink.ready
			sink_channel       => id_router_004_src_channel,             --          .channel
			sink_data          => id_router_004_src_data,                --          .data
			sink_startofpacket => id_router_004_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_004_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_004_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_004_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_004_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_004_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_004_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_004_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_004_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_004_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_004_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_004_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_004_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_004_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_004_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_005 : component p2_grms_qsys_rsp_xbar_demux
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_005_src_ready,               --      sink.ready
			sink_channel       => id_router_005_src_channel,             --          .channel
			sink_data          => id_router_005_src_data,                --          .data
			sink_startofpacket => id_router_005_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_005_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_005_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_005_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_005_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_005_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_005_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_005_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_005_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_005_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_005_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_005_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_005_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_005_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_005_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_006 : component p2_grms_qsys_rsp_xbar_demux
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_006_src_ready,               --      sink.ready
			sink_channel       => id_router_006_src_channel,             --          .channel
			sink_data          => id_router_006_src_data,                --          .data
			sink_startofpacket => id_router_006_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_006_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_006_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_006_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_006_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_006_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_006_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_006_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_006_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_006_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_006_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_006_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_006_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_006_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_006_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_007 : component p2_grms_qsys_rsp_xbar_demux
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_007_src_ready,               --      sink.ready
			sink_channel       => id_router_007_src_channel,             --          .channel
			sink_data          => id_router_007_src_data,                --          .data
			sink_startofpacket => id_router_007_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_007_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_007_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_007_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_007_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_007_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_007_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_007_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_007_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_007_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_007_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_007_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_007_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_007_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_007_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_008 : component p2_grms_qsys_rsp_xbar_demux
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_008_src_ready,               --      sink.ready
			sink_channel       => id_router_008_src_channel,             --          .channel
			sink_data          => id_router_008_src_data,                --          .data
			sink_startofpacket => id_router_008_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_008_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_008_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_008_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_008_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_008_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_008_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_008_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_008_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_008_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_008_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_008_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_008_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_008_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_008_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_009 : component p2_grms_qsys_rsp_xbar_demux
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_009_src_ready,               --      sink.ready
			sink_channel       => id_router_009_src_channel,             --          .channel
			sink_data          => id_router_009_src_data,                --          .data
			sink_startofpacket => id_router_009_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_009_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_009_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_009_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_009_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_009_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_009_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_009_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_009_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_009_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_009_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_009_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_009_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_009_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_009_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_010 : component p2_grms_qsys_rsp_xbar_demux
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_010_src_ready,               --      sink.ready
			sink_channel       => id_router_010_src_channel,             --          .channel
			sink_data          => id_router_010_src_data,                --          .data
			sink_startofpacket => id_router_010_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_010_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_010_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_010_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_010_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_010_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_010_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_010_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_010_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_010_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_010_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_010_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_010_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_010_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_010_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_011 : component p2_grms_qsys_rsp_xbar_demux
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_011_src_ready,               --      sink.ready
			sink_channel       => id_router_011_src_channel,             --          .channel
			sink_data          => id_router_011_src_data,                --          .data
			sink_startofpacket => id_router_011_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_011_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_011_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_011_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_011_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_011_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_011_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_011_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_011_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_011_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_011_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_011_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_011_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_011_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_011_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_012 : component p2_grms_qsys_rsp_xbar_demux
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_012_src_ready,               --      sink.ready
			sink_channel       => id_router_012_src_channel,             --          .channel
			sink_data          => id_router_012_src_data,                --          .data
			sink_startofpacket => id_router_012_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_012_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_012_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_012_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_012_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_012_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_012_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_012_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_012_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_012_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_012_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_012_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_012_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_012_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_012_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_013 : component p2_grms_qsys_rsp_xbar_demux
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_013_src_ready,               --      sink.ready
			sink_channel       => id_router_013_src_channel,             --          .channel
			sink_data          => id_router_013_src_data,                --          .data
			sink_startofpacket => id_router_013_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_013_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_013_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_013_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_013_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_013_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_013_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_013_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_013_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_013_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_013_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_013_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_013_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_013_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_013_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_mux : component p2_grms_qsys_rsp_xbar_mux
		port map (
			clk                  => clk_clk,                               --       clk.clk
			reset                => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready            => rsp_xbar_mux_src_ready,                --       src.ready
			src_valid            => rsp_xbar_mux_src_valid,                --          .valid
			src_data             => rsp_xbar_mux_src_data,                 --          .data
			src_channel          => rsp_xbar_mux_src_channel,              --          .channel
			src_startofpacket    => rsp_xbar_mux_src_startofpacket,        --          .startofpacket
			src_endofpacket      => rsp_xbar_mux_src_endofpacket,          --          .endofpacket
			sink0_ready          => rsp_xbar_demux_src0_ready,             --     sink0.ready
			sink0_valid          => rsp_xbar_demux_src0_valid,             --          .valid
			sink0_channel        => rsp_xbar_demux_src0_channel,           --          .channel
			sink0_data           => rsp_xbar_demux_src0_data,              --          .data
			sink0_startofpacket  => rsp_xbar_demux_src0_startofpacket,     --          .startofpacket
			sink0_endofpacket    => rsp_xbar_demux_src0_endofpacket,       --          .endofpacket
			sink1_ready          => rsp_xbar_demux_001_src0_ready,         --     sink1.ready
			sink1_valid          => rsp_xbar_demux_001_src0_valid,         --          .valid
			sink1_channel        => rsp_xbar_demux_001_src0_channel,       --          .channel
			sink1_data           => rsp_xbar_demux_001_src0_data,          --          .data
			sink1_startofpacket  => rsp_xbar_demux_001_src0_startofpacket, --          .startofpacket
			sink1_endofpacket    => rsp_xbar_demux_001_src0_endofpacket,   --          .endofpacket
			sink2_ready          => rsp_xbar_demux_002_src0_ready,         --     sink2.ready
			sink2_valid          => rsp_xbar_demux_002_src0_valid,         --          .valid
			sink2_channel        => rsp_xbar_demux_002_src0_channel,       --          .channel
			sink2_data           => rsp_xbar_demux_002_src0_data,          --          .data
			sink2_startofpacket  => rsp_xbar_demux_002_src0_startofpacket, --          .startofpacket
			sink2_endofpacket    => rsp_xbar_demux_002_src0_endofpacket,   --          .endofpacket
			sink3_ready          => rsp_xbar_demux_003_src0_ready,         --     sink3.ready
			sink3_valid          => rsp_xbar_demux_003_src0_valid,         --          .valid
			sink3_channel        => rsp_xbar_demux_003_src0_channel,       --          .channel
			sink3_data           => rsp_xbar_demux_003_src0_data,          --          .data
			sink3_startofpacket  => rsp_xbar_demux_003_src0_startofpacket, --          .startofpacket
			sink3_endofpacket    => rsp_xbar_demux_003_src0_endofpacket,   --          .endofpacket
			sink4_ready          => rsp_xbar_demux_004_src0_ready,         --     sink4.ready
			sink4_valid          => rsp_xbar_demux_004_src0_valid,         --          .valid
			sink4_channel        => rsp_xbar_demux_004_src0_channel,       --          .channel
			sink4_data           => rsp_xbar_demux_004_src0_data,          --          .data
			sink4_startofpacket  => rsp_xbar_demux_004_src0_startofpacket, --          .startofpacket
			sink4_endofpacket    => rsp_xbar_demux_004_src0_endofpacket,   --          .endofpacket
			sink5_ready          => rsp_xbar_demux_005_src0_ready,         --     sink5.ready
			sink5_valid          => rsp_xbar_demux_005_src0_valid,         --          .valid
			sink5_channel        => rsp_xbar_demux_005_src0_channel,       --          .channel
			sink5_data           => rsp_xbar_demux_005_src0_data,          --          .data
			sink5_startofpacket  => rsp_xbar_demux_005_src0_startofpacket, --          .startofpacket
			sink5_endofpacket    => rsp_xbar_demux_005_src0_endofpacket,   --          .endofpacket
			sink6_ready          => rsp_xbar_demux_006_src0_ready,         --     sink6.ready
			sink6_valid          => rsp_xbar_demux_006_src0_valid,         --          .valid
			sink6_channel        => rsp_xbar_demux_006_src0_channel,       --          .channel
			sink6_data           => rsp_xbar_demux_006_src0_data,          --          .data
			sink6_startofpacket  => rsp_xbar_demux_006_src0_startofpacket, --          .startofpacket
			sink6_endofpacket    => rsp_xbar_demux_006_src0_endofpacket,   --          .endofpacket
			sink7_ready          => rsp_xbar_demux_007_src0_ready,         --     sink7.ready
			sink7_valid          => rsp_xbar_demux_007_src0_valid,         --          .valid
			sink7_channel        => rsp_xbar_demux_007_src0_channel,       --          .channel
			sink7_data           => rsp_xbar_demux_007_src0_data,          --          .data
			sink7_startofpacket  => rsp_xbar_demux_007_src0_startofpacket, --          .startofpacket
			sink7_endofpacket    => rsp_xbar_demux_007_src0_endofpacket,   --          .endofpacket
			sink8_ready          => rsp_xbar_demux_008_src0_ready,         --     sink8.ready
			sink8_valid          => rsp_xbar_demux_008_src0_valid,         --          .valid
			sink8_channel        => rsp_xbar_demux_008_src0_channel,       --          .channel
			sink8_data           => rsp_xbar_demux_008_src0_data,          --          .data
			sink8_startofpacket  => rsp_xbar_demux_008_src0_startofpacket, --          .startofpacket
			sink8_endofpacket    => rsp_xbar_demux_008_src0_endofpacket,   --          .endofpacket
			sink9_ready          => rsp_xbar_demux_009_src0_ready,         --     sink9.ready
			sink9_valid          => rsp_xbar_demux_009_src0_valid,         --          .valid
			sink9_channel        => rsp_xbar_demux_009_src0_channel,       --          .channel
			sink9_data           => rsp_xbar_demux_009_src0_data,          --          .data
			sink9_startofpacket  => rsp_xbar_demux_009_src0_startofpacket, --          .startofpacket
			sink9_endofpacket    => rsp_xbar_demux_009_src0_endofpacket,   --          .endofpacket
			sink10_ready         => rsp_xbar_demux_010_src0_ready,         --    sink10.ready
			sink10_valid         => rsp_xbar_demux_010_src0_valid,         --          .valid
			sink10_channel       => rsp_xbar_demux_010_src0_channel,       --          .channel
			sink10_data          => rsp_xbar_demux_010_src0_data,          --          .data
			sink10_startofpacket => rsp_xbar_demux_010_src0_startofpacket, --          .startofpacket
			sink10_endofpacket   => rsp_xbar_demux_010_src0_endofpacket,   --          .endofpacket
			sink11_ready         => rsp_xbar_demux_011_src0_ready,         --    sink11.ready
			sink11_valid         => rsp_xbar_demux_011_src0_valid,         --          .valid
			sink11_channel       => rsp_xbar_demux_011_src0_channel,       --          .channel
			sink11_data          => rsp_xbar_demux_011_src0_data,          --          .data
			sink11_startofpacket => rsp_xbar_demux_011_src0_startofpacket, --          .startofpacket
			sink11_endofpacket   => rsp_xbar_demux_011_src0_endofpacket,   --          .endofpacket
			sink12_ready         => rsp_xbar_demux_012_src0_ready,         --    sink12.ready
			sink12_valid         => rsp_xbar_demux_012_src0_valid,         --          .valid
			sink12_channel       => rsp_xbar_demux_012_src0_channel,       --          .channel
			sink12_data          => rsp_xbar_demux_012_src0_data,          --          .data
			sink12_startofpacket => rsp_xbar_demux_012_src0_startofpacket, --          .startofpacket
			sink12_endofpacket   => rsp_xbar_demux_012_src0_endofpacket,   --          .endofpacket
			sink13_ready         => rsp_xbar_demux_013_src0_ready,         --    sink13.ready
			sink13_valid         => rsp_xbar_demux_013_src0_valid,         --          .valid
			sink13_channel       => rsp_xbar_demux_013_src0_channel,       --          .channel
			sink13_data          => rsp_xbar_demux_013_src0_data,          --          .data
			sink13_startofpacket => rsp_xbar_demux_013_src0_startofpacket, --          .startofpacket
			sink13_endofpacket   => rsp_xbar_demux_013_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_mux_001 : component p2_grms_qsys_rsp_xbar_mux
		port map (
			clk                  => clk_clk,                               --       clk.clk
			reset                => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready            => rsp_xbar_mux_001_src_ready,            --       src.ready
			src_valid            => rsp_xbar_mux_001_src_valid,            --          .valid
			src_data             => rsp_xbar_mux_001_src_data,             --          .data
			src_channel          => rsp_xbar_mux_001_src_channel,          --          .channel
			src_startofpacket    => rsp_xbar_mux_001_src_startofpacket,    --          .startofpacket
			src_endofpacket      => rsp_xbar_mux_001_src_endofpacket,      --          .endofpacket
			sink0_ready          => rsp_xbar_demux_src1_ready,             --     sink0.ready
			sink0_valid          => rsp_xbar_demux_src1_valid,             --          .valid
			sink0_channel        => rsp_xbar_demux_src1_channel,           --          .channel
			sink0_data           => rsp_xbar_demux_src1_data,              --          .data
			sink0_startofpacket  => rsp_xbar_demux_src1_startofpacket,     --          .startofpacket
			sink0_endofpacket    => rsp_xbar_demux_src1_endofpacket,       --          .endofpacket
			sink1_ready          => rsp_xbar_demux_001_src1_ready,         --     sink1.ready
			sink1_valid          => rsp_xbar_demux_001_src1_valid,         --          .valid
			sink1_channel        => rsp_xbar_demux_001_src1_channel,       --          .channel
			sink1_data           => rsp_xbar_demux_001_src1_data,          --          .data
			sink1_startofpacket  => rsp_xbar_demux_001_src1_startofpacket, --          .startofpacket
			sink1_endofpacket    => rsp_xbar_demux_001_src1_endofpacket,   --          .endofpacket
			sink2_ready          => rsp_xbar_demux_002_src1_ready,         --     sink2.ready
			sink2_valid          => rsp_xbar_demux_002_src1_valid,         --          .valid
			sink2_channel        => rsp_xbar_demux_002_src1_channel,       --          .channel
			sink2_data           => rsp_xbar_demux_002_src1_data,          --          .data
			sink2_startofpacket  => rsp_xbar_demux_002_src1_startofpacket, --          .startofpacket
			sink2_endofpacket    => rsp_xbar_demux_002_src1_endofpacket,   --          .endofpacket
			sink3_ready          => rsp_xbar_demux_003_src1_ready,         --     sink3.ready
			sink3_valid          => rsp_xbar_demux_003_src1_valid,         --          .valid
			sink3_channel        => rsp_xbar_demux_003_src1_channel,       --          .channel
			sink3_data           => rsp_xbar_demux_003_src1_data,          --          .data
			sink3_startofpacket  => rsp_xbar_demux_003_src1_startofpacket, --          .startofpacket
			sink3_endofpacket    => rsp_xbar_demux_003_src1_endofpacket,   --          .endofpacket
			sink4_ready          => rsp_xbar_demux_004_src1_ready,         --     sink4.ready
			sink4_valid          => rsp_xbar_demux_004_src1_valid,         --          .valid
			sink4_channel        => rsp_xbar_demux_004_src1_channel,       --          .channel
			sink4_data           => rsp_xbar_demux_004_src1_data,          --          .data
			sink4_startofpacket  => rsp_xbar_demux_004_src1_startofpacket, --          .startofpacket
			sink4_endofpacket    => rsp_xbar_demux_004_src1_endofpacket,   --          .endofpacket
			sink5_ready          => rsp_xbar_demux_005_src1_ready,         --     sink5.ready
			sink5_valid          => rsp_xbar_demux_005_src1_valid,         --          .valid
			sink5_channel        => rsp_xbar_demux_005_src1_channel,       --          .channel
			sink5_data           => rsp_xbar_demux_005_src1_data,          --          .data
			sink5_startofpacket  => rsp_xbar_demux_005_src1_startofpacket, --          .startofpacket
			sink5_endofpacket    => rsp_xbar_demux_005_src1_endofpacket,   --          .endofpacket
			sink6_ready          => rsp_xbar_demux_006_src1_ready,         --     sink6.ready
			sink6_valid          => rsp_xbar_demux_006_src1_valid,         --          .valid
			sink6_channel        => rsp_xbar_demux_006_src1_channel,       --          .channel
			sink6_data           => rsp_xbar_demux_006_src1_data,          --          .data
			sink6_startofpacket  => rsp_xbar_demux_006_src1_startofpacket, --          .startofpacket
			sink6_endofpacket    => rsp_xbar_demux_006_src1_endofpacket,   --          .endofpacket
			sink7_ready          => rsp_xbar_demux_007_src1_ready,         --     sink7.ready
			sink7_valid          => rsp_xbar_demux_007_src1_valid,         --          .valid
			sink7_channel        => rsp_xbar_demux_007_src1_channel,       --          .channel
			sink7_data           => rsp_xbar_demux_007_src1_data,          --          .data
			sink7_startofpacket  => rsp_xbar_demux_007_src1_startofpacket, --          .startofpacket
			sink7_endofpacket    => rsp_xbar_demux_007_src1_endofpacket,   --          .endofpacket
			sink8_ready          => rsp_xbar_demux_008_src1_ready,         --     sink8.ready
			sink8_valid          => rsp_xbar_demux_008_src1_valid,         --          .valid
			sink8_channel        => rsp_xbar_demux_008_src1_channel,       --          .channel
			sink8_data           => rsp_xbar_demux_008_src1_data,          --          .data
			sink8_startofpacket  => rsp_xbar_demux_008_src1_startofpacket, --          .startofpacket
			sink8_endofpacket    => rsp_xbar_demux_008_src1_endofpacket,   --          .endofpacket
			sink9_ready          => rsp_xbar_demux_009_src1_ready,         --     sink9.ready
			sink9_valid          => rsp_xbar_demux_009_src1_valid,         --          .valid
			sink9_channel        => rsp_xbar_demux_009_src1_channel,       --          .channel
			sink9_data           => rsp_xbar_demux_009_src1_data,          --          .data
			sink9_startofpacket  => rsp_xbar_demux_009_src1_startofpacket, --          .startofpacket
			sink9_endofpacket    => rsp_xbar_demux_009_src1_endofpacket,   --          .endofpacket
			sink10_ready         => rsp_xbar_demux_010_src1_ready,         --    sink10.ready
			sink10_valid         => rsp_xbar_demux_010_src1_valid,         --          .valid
			sink10_channel       => rsp_xbar_demux_010_src1_channel,       --          .channel
			sink10_data          => rsp_xbar_demux_010_src1_data,          --          .data
			sink10_startofpacket => rsp_xbar_demux_010_src1_startofpacket, --          .startofpacket
			sink10_endofpacket   => rsp_xbar_demux_010_src1_endofpacket,   --          .endofpacket
			sink11_ready         => rsp_xbar_demux_011_src1_ready,         --    sink11.ready
			sink11_valid         => rsp_xbar_demux_011_src1_valid,         --          .valid
			sink11_channel       => rsp_xbar_demux_011_src1_channel,       --          .channel
			sink11_data          => rsp_xbar_demux_011_src1_data,          --          .data
			sink11_startofpacket => rsp_xbar_demux_011_src1_startofpacket, --          .startofpacket
			sink11_endofpacket   => rsp_xbar_demux_011_src1_endofpacket,   --          .endofpacket
			sink12_ready         => rsp_xbar_demux_012_src1_ready,         --    sink12.ready
			sink12_valid         => rsp_xbar_demux_012_src1_valid,         --          .valid
			sink12_channel       => rsp_xbar_demux_012_src1_channel,       --          .channel
			sink12_data          => rsp_xbar_demux_012_src1_data,          --          .data
			sink12_startofpacket => rsp_xbar_demux_012_src1_startofpacket, --          .startofpacket
			sink12_endofpacket   => rsp_xbar_demux_012_src1_endofpacket,   --          .endofpacket
			sink13_ready         => rsp_xbar_demux_013_src1_ready,         --    sink13.ready
			sink13_valid         => rsp_xbar_demux_013_src1_valid,         --          .valid
			sink13_channel       => rsp_xbar_demux_013_src1_channel,       --          .channel
			sink13_data          => rsp_xbar_demux_013_src1_data,          --          .data
			sink13_startofpacket => rsp_xbar_demux_013_src1_startofpacket, --          .startofpacket
			sink13_endofpacket   => rsp_xbar_demux_013_src1_endofpacket    --          .endofpacket
		);

	width_adapter : component p2_grms_qsys_width_adapter
		generic map (
			IN_PKT_ADDR_H                 => 60,
			IN_PKT_ADDR_L                 => 36,
			IN_PKT_DATA_H                 => 31,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 35,
			IN_PKT_BYTEEN_L               => 32,
			IN_PKT_BYTE_CNT_H             => 69,
			IN_PKT_BYTE_CNT_L             => 67,
			IN_PKT_TRANS_COMPRESSED_READ  => 61,
			IN_PKT_BURSTWRAP_H            => 72,
			IN_PKT_BURSTWRAP_L            => 70,
			IN_PKT_BURST_SIZE_H           => 75,
			IN_PKT_BURST_SIZE_L           => 73,
			IN_PKT_RESPONSE_STATUS_H      => 99,
			IN_PKT_RESPONSE_STATUS_L      => 98,
			IN_PKT_TRANS_EXCLUSIVE        => 66,
			IN_PKT_BURST_TYPE_H           => 77,
			IN_PKT_BURST_TYPE_L           => 76,
			IN_ST_DATA_W                  => 100,
			OUT_PKT_ADDR_H                => 42,
			OUT_PKT_ADDR_L                => 18,
			OUT_PKT_DATA_H                => 15,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 17,
			OUT_PKT_BYTEEN_L              => 16,
			OUT_PKT_BYTE_CNT_H            => 51,
			OUT_PKT_BYTE_CNT_L            => 49,
			OUT_PKT_TRANS_COMPRESSED_READ => 43,
			OUT_PKT_BURST_SIZE_H          => 57,
			OUT_PKT_BURST_SIZE_L          => 55,
			OUT_PKT_RESPONSE_STATUS_H     => 81,
			OUT_PKT_RESPONSE_STATUS_L     => 80,
			OUT_PKT_TRANS_EXCLUSIVE       => 48,
			OUT_PKT_BURST_TYPE_H          => 59,
			OUT_PKT_BURST_TYPE_L          => 58,
			OUT_ST_DATA_W                 => 82,
			ST_CHANNEL_W                  => 14,
			OPTIMIZE_FOR_RSP              => 0,
			RESPONSE_PATH                 => 0
		)
		port map (
			clk                  => clk_clk,                            --       clk.clk
			reset                => rst_controller_reset_out_reset,     -- clk_reset.reset
			in_valid             => cmd_xbar_mux_002_src_valid,         --      sink.valid
			in_channel           => cmd_xbar_mux_002_src_channel,       --          .channel
			in_startofpacket     => cmd_xbar_mux_002_src_startofpacket, --          .startofpacket
			in_endofpacket       => cmd_xbar_mux_002_src_endofpacket,   --          .endofpacket
			in_ready             => cmd_xbar_mux_002_src_ready,         --          .ready
			in_data              => cmd_xbar_mux_002_src_data,          --          .data
			out_endofpacket      => width_adapter_src_endofpacket,      --       src.endofpacket
			out_data             => width_adapter_src_data,             --          .data
			out_channel          => width_adapter_src_channel,          --          .channel
			out_valid            => width_adapter_src_valid,            --          .valid
			out_ready            => width_adapter_src_ready,            --          .ready
			out_startofpacket    => width_adapter_src_startofpacket,    --          .startofpacket
			in_command_size_data => "000"                               -- (terminated)
		);

	width_adapter_001 : component p2_grms_qsys_width_adapter_001
		generic map (
			IN_PKT_ADDR_H                 => 42,
			IN_PKT_ADDR_L                 => 18,
			IN_PKT_DATA_H                 => 15,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 17,
			IN_PKT_BYTEEN_L               => 16,
			IN_PKT_BYTE_CNT_H             => 51,
			IN_PKT_BYTE_CNT_L             => 49,
			IN_PKT_TRANS_COMPRESSED_READ  => 43,
			IN_PKT_BURSTWRAP_H            => 54,
			IN_PKT_BURSTWRAP_L            => 52,
			IN_PKT_BURST_SIZE_H           => 57,
			IN_PKT_BURST_SIZE_L           => 55,
			IN_PKT_RESPONSE_STATUS_H      => 81,
			IN_PKT_RESPONSE_STATUS_L      => 80,
			IN_PKT_TRANS_EXCLUSIVE        => 48,
			IN_PKT_BURST_TYPE_H           => 59,
			IN_PKT_BURST_TYPE_L           => 58,
			IN_ST_DATA_W                  => 82,
			OUT_PKT_ADDR_H                => 60,
			OUT_PKT_ADDR_L                => 36,
			OUT_PKT_DATA_H                => 31,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 35,
			OUT_PKT_BYTEEN_L              => 32,
			OUT_PKT_BYTE_CNT_H            => 69,
			OUT_PKT_BYTE_CNT_L            => 67,
			OUT_PKT_TRANS_COMPRESSED_READ => 61,
			OUT_PKT_BURST_SIZE_H          => 75,
			OUT_PKT_BURST_SIZE_L          => 73,
			OUT_PKT_RESPONSE_STATUS_H     => 99,
			OUT_PKT_RESPONSE_STATUS_L     => 98,
			OUT_PKT_TRANS_EXCLUSIVE       => 66,
			OUT_PKT_BURST_TYPE_H          => 77,
			OUT_PKT_BURST_TYPE_L          => 76,
			OUT_ST_DATA_W                 => 100,
			ST_CHANNEL_W                  => 14,
			OPTIMIZE_FOR_RSP              => 1,
			RESPONSE_PATH                 => 1
		)
		port map (
			clk                  => clk_clk,                             --       clk.clk
			reset                => rst_controller_reset_out_reset,      -- clk_reset.reset
			in_valid             => id_router_002_src_valid,             --      sink.valid
			in_channel           => id_router_002_src_channel,           --          .channel
			in_startofpacket     => id_router_002_src_startofpacket,     --          .startofpacket
			in_endofpacket       => id_router_002_src_endofpacket,       --          .endofpacket
			in_ready             => id_router_002_src_ready,             --          .ready
			in_data              => id_router_002_src_data,              --          .data
			out_endofpacket      => width_adapter_001_src_endofpacket,   --       src.endofpacket
			out_data             => width_adapter_001_src_data,          --          .data
			out_channel          => width_adapter_001_src_channel,       --          .channel
			out_valid            => width_adapter_001_src_valid,         --          .valid
			out_ready            => width_adapter_001_src_ready,         --          .ready
			out_startofpacket    => width_adapter_001_src_startofpacket, --          .startofpacket
			in_command_size_data => "000"                                -- (terminated)
		);

	irq_mapper : component p2_grms_qsys_irq_mapper
		port map (
			clk           => clk_clk,                        --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			sender_irq    => nios2_qsys_grms_d_irq_irq       --    sender.irq
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	jtag_uart_grms_avalon_jtag_slave_translator_avalon_anti_slave_0_write_ports_inv <= not jtag_uart_grms_avalon_jtag_slave_translator_avalon_anti_slave_0_write;

	jtag_uart_grms_avalon_jtag_slave_translator_avalon_anti_slave_0_read_ports_inv <= not jtag_uart_grms_avalon_jtag_slave_translator_avalon_anti_slave_0_read;

	new_sdram_controller_grms_s1_translator_avalon_anti_slave_0_write_ports_inv <= not new_sdram_controller_grms_s1_translator_avalon_anti_slave_0_write;

	new_sdram_controller_grms_s1_translator_avalon_anti_slave_0_read_ports_inv <= not new_sdram_controller_grms_s1_translator_avalon_anti_slave_0_read;

	new_sdram_controller_grms_s1_translator_avalon_anti_slave_0_byteenable_ports_inv <= not new_sdram_controller_grms_s1_translator_avalon_anti_slave_0_byteenable;

	timer_grms_s1_translator_avalon_anti_slave_0_write_ports_inv <= not timer_grms_s1_translator_avalon_anti_slave_0_write;

	pc_grms_s1_translator_avalon_anti_slave_0_write_ports_inv <= not pc_grms_s1_translator_avalon_anti_slave_0_write;

	pd_grms_s1_translator_avalon_anti_slave_0_write_ports_inv <= not pd_grms_s1_translator_avalon_anti_slave_0_write;

	pe_grms_s1_translator_avalon_anti_slave_0_write_ports_inv <= not pe_grms_s1_translator_avalon_anti_slave_0_write;

	pf_grms_s1_translator_avalon_anti_slave_0_write_ports_inv <= not pf_grms_s1_translator_avalon_anti_slave_0_write;

	pg_grms_s1_translator_avalon_anti_slave_0_write_ports_inv <= not pg_grms_s1_translator_avalon_anti_slave_0_write;

	ph_grms_s1_translator_avalon_anti_slave_0_write_ports_inv <= not ph_grms_s1_translator_avalon_anti_slave_0_write;

	pi_grms_s1_translator_avalon_anti_slave_0_write_ports_inv <= not pi_grms_s1_translator_avalon_anti_slave_0_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of p2_grms_qsys
